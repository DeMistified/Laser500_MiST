
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"00",x"00",x"00",x"40"),
     1 => (x"fd",x"80",x"80",x"80"),
     2 => (x"00",x"00",x"00",x"7d"),
     3 => (x"38",x"10",x"7f",x"7f"),
     4 => (x"00",x"00",x"44",x"6c"),
     5 => (x"7f",x"3f",x"00",x"00"),
     6 => (x"7c",x"00",x"00",x"40"),
     7 => (x"0c",x"18",x"0c",x"7c"),
     8 => (x"00",x"00",x"78",x"7c"),
     9 => (x"04",x"04",x"7c",x"7c"),
    10 => (x"00",x"00",x"78",x"7c"),
    11 => (x"44",x"44",x"7c",x"38"),
    12 => (x"00",x"00",x"38",x"7c"),
    13 => (x"24",x"24",x"fc",x"fc"),
    14 => (x"00",x"00",x"18",x"3c"),
    15 => (x"24",x"24",x"3c",x"18"),
    16 => (x"00",x"00",x"fc",x"fc"),
    17 => (x"04",x"04",x"7c",x"7c"),
    18 => (x"00",x"00",x"08",x"0c"),
    19 => (x"54",x"54",x"5c",x"48"),
    20 => (x"00",x"00",x"20",x"74"),
    21 => (x"44",x"7f",x"3f",x"04"),
    22 => (x"00",x"00",x"00",x"44"),
    23 => (x"40",x"40",x"7c",x"3c"),
    24 => (x"00",x"00",x"7c",x"7c"),
    25 => (x"60",x"60",x"3c",x"1c"),
    26 => (x"3c",x"00",x"1c",x"3c"),
    27 => (x"60",x"30",x"60",x"7c"),
    28 => (x"44",x"00",x"3c",x"7c"),
    29 => (x"38",x"10",x"38",x"6c"),
    30 => (x"00",x"00",x"44",x"6c"),
    31 => (x"60",x"e0",x"bc",x"1c"),
    32 => (x"00",x"00",x"1c",x"3c"),
    33 => (x"5c",x"74",x"64",x"44"),
    34 => (x"00",x"00",x"44",x"4c"),
    35 => (x"77",x"3e",x"08",x"08"),
    36 => (x"00",x"00",x"41",x"41"),
    37 => (x"7f",x"7f",x"00",x"00"),
    38 => (x"00",x"00",x"00",x"00"),
    39 => (x"3e",x"77",x"41",x"41"),
    40 => (x"02",x"00",x"08",x"08"),
    41 => (x"02",x"03",x"01",x"01"),
    42 => (x"7f",x"00",x"01",x"02"),
    43 => (x"7f",x"7f",x"7f",x"7f"),
    44 => (x"08",x"00",x"7f",x"7f"),
    45 => (x"3e",x"1c",x"1c",x"08"),
    46 => (x"7f",x"7f",x"7f",x"3e"),
    47 => (x"1c",x"3e",x"3e",x"7f"),
    48 => (x"00",x"08",x"08",x"1c"),
    49 => (x"7c",x"7c",x"18",x"10"),
    50 => (x"00",x"00",x"10",x"18"),
    51 => (x"7c",x"7c",x"30",x"10"),
    52 => (x"10",x"00",x"10",x"30"),
    53 => (x"78",x"60",x"60",x"30"),
    54 => (x"42",x"00",x"06",x"1e"),
    55 => (x"3c",x"18",x"3c",x"66"),
    56 => (x"78",x"00",x"42",x"66"),
    57 => (x"c6",x"c2",x"6a",x"38"),
    58 => (x"60",x"00",x"38",x"6c"),
    59 => (x"00",x"60",x"00",x"00"),
    60 => (x"0e",x"00",x"60",x"00"),
    61 => (x"5d",x"5c",x"5b",x"5e"),
    62 => (x"4c",x"71",x"1e",x"0e"),
    63 => (x"bf",x"ed",x"ed",x"c2"),
    64 => (x"c0",x"4b",x"c0",x"4d"),
    65 => (x"02",x"ab",x"74",x"1e"),
    66 => (x"a6",x"c4",x"87",x"c7"),
    67 => (x"c5",x"78",x"c0",x"48"),
    68 => (x"48",x"a6",x"c4",x"87"),
    69 => (x"66",x"c4",x"78",x"c1"),
    70 => (x"ee",x"49",x"73",x"1e"),
    71 => (x"86",x"c8",x"87",x"df"),
    72 => (x"ef",x"49",x"e0",x"c0"),
    73 => (x"a5",x"c4",x"87",x"ef"),
    74 => (x"f0",x"49",x"6a",x"4a"),
    75 => (x"c6",x"f1",x"87",x"f0"),
    76 => (x"c1",x"85",x"cb",x"87"),
    77 => (x"ab",x"b7",x"c8",x"83"),
    78 => (x"87",x"c7",x"ff",x"04"),
    79 => (x"26",x"4d",x"26",x"26"),
    80 => (x"26",x"4b",x"26",x"4c"),
    81 => (x"4a",x"71",x"1e",x"4f"),
    82 => (x"5a",x"f1",x"ed",x"c2"),
    83 => (x"48",x"f1",x"ed",x"c2"),
    84 => (x"fe",x"49",x"78",x"c7"),
    85 => (x"4f",x"26",x"87",x"dd"),
    86 => (x"71",x"1e",x"73",x"1e"),
    87 => (x"aa",x"b7",x"c0",x"4a"),
    88 => (x"c2",x"87",x"d3",x"03"),
    89 => (x"05",x"bf",x"e8",x"d2"),
    90 => (x"4b",x"c1",x"87",x"c4"),
    91 => (x"4b",x"c0",x"87",x"c2"),
    92 => (x"5b",x"ec",x"d2",x"c2"),
    93 => (x"d2",x"c2",x"87",x"c4"),
    94 => (x"d2",x"c2",x"5a",x"ec"),
    95 => (x"c1",x"4a",x"bf",x"e8"),
    96 => (x"a2",x"c0",x"c1",x"9a"),
    97 => (x"87",x"e8",x"ec",x"49"),
    98 => (x"d2",x"c2",x"48",x"fc"),
    99 => (x"fe",x"78",x"bf",x"e8"),
   100 => (x"71",x"1e",x"87",x"ef"),
   101 => (x"1e",x"66",x"c4",x"4a"),
   102 => (x"f9",x"e9",x"49",x"72"),
   103 => (x"4f",x"26",x"26",x"87"),
   104 => (x"e8",x"d2",x"c2",x"1e"),
   105 => (x"db",x"e6",x"49",x"bf"),
   106 => (x"e5",x"ed",x"c2",x"87"),
   107 => (x"78",x"bf",x"e8",x"48"),
   108 => (x"48",x"e1",x"ed",x"c2"),
   109 => (x"c2",x"78",x"bf",x"ec"),
   110 => (x"4a",x"bf",x"e5",x"ed"),
   111 => (x"99",x"ff",x"c3",x"49"),
   112 => (x"72",x"2a",x"b7",x"c8"),
   113 => (x"c2",x"b0",x"71",x"48"),
   114 => (x"26",x"58",x"ed",x"ed"),
   115 => (x"5b",x"5e",x"0e",x"4f"),
   116 => (x"71",x"0e",x"5d",x"5c"),
   117 => (x"87",x"c8",x"ff",x"4b"),
   118 => (x"48",x"e0",x"ed",x"c2"),
   119 => (x"49",x"73",x"50",x"c0"),
   120 => (x"70",x"87",x"c1",x"e6"),
   121 => (x"9c",x"c2",x"4c",x"49"),
   122 => (x"cb",x"49",x"ee",x"cb"),
   123 => (x"49",x"70",x"87",x"c2"),
   124 => (x"e0",x"ed",x"c2",x"4d"),
   125 => (x"c1",x"05",x"bf",x"97"),
   126 => (x"66",x"d0",x"87",x"e2"),
   127 => (x"e9",x"ed",x"c2",x"49"),
   128 => (x"d6",x"05",x"99",x"bf"),
   129 => (x"49",x"66",x"d4",x"87"),
   130 => (x"bf",x"e1",x"ed",x"c2"),
   131 => (x"87",x"cb",x"05",x"99"),
   132 => (x"cf",x"e5",x"49",x"73"),
   133 => (x"02",x"98",x"70",x"87"),
   134 => (x"c1",x"87",x"c1",x"c1"),
   135 => (x"87",x"c0",x"fe",x"4c"),
   136 => (x"d7",x"ca",x"49",x"75"),
   137 => (x"02",x"98",x"70",x"87"),
   138 => (x"ed",x"c2",x"87",x"c6"),
   139 => (x"50",x"c1",x"48",x"e0"),
   140 => (x"97",x"e0",x"ed",x"c2"),
   141 => (x"e3",x"c0",x"05",x"bf"),
   142 => (x"e9",x"ed",x"c2",x"87"),
   143 => (x"66",x"d0",x"49",x"bf"),
   144 => (x"d6",x"ff",x"05",x"99"),
   145 => (x"e1",x"ed",x"c2",x"87"),
   146 => (x"66",x"d4",x"49",x"bf"),
   147 => (x"ca",x"ff",x"05",x"99"),
   148 => (x"e4",x"49",x"73",x"87"),
   149 => (x"98",x"70",x"87",x"ce"),
   150 => (x"87",x"ff",x"fe",x"05"),
   151 => (x"dc",x"fb",x"48",x"74"),
   152 => (x"5b",x"5e",x"0e",x"87"),
   153 => (x"f4",x"0e",x"5d",x"5c"),
   154 => (x"4c",x"4d",x"c0",x"86"),
   155 => (x"c4",x"7e",x"bf",x"ec"),
   156 => (x"ed",x"c2",x"48",x"a6"),
   157 => (x"c1",x"78",x"bf",x"ed"),
   158 => (x"c7",x"1e",x"c0",x"1e"),
   159 => (x"87",x"cd",x"fd",x"49"),
   160 => (x"98",x"70",x"86",x"c8"),
   161 => (x"ff",x"87",x"cd",x"02"),
   162 => (x"87",x"cc",x"fb",x"49"),
   163 => (x"e3",x"49",x"da",x"c1"),
   164 => (x"4d",x"c1",x"87",x"d2"),
   165 => (x"97",x"e0",x"ed",x"c2"),
   166 => (x"87",x"c3",x"02",x"bf"),
   167 => (x"c2",x"87",x"fb",x"cf"),
   168 => (x"4b",x"bf",x"e5",x"ed"),
   169 => (x"bf",x"e8",x"d2",x"c2"),
   170 => (x"87",x"e9",x"c0",x"05"),
   171 => (x"e2",x"49",x"fd",x"c3"),
   172 => (x"fa",x"c3",x"87",x"f2"),
   173 => (x"87",x"ec",x"e2",x"49"),
   174 => (x"ff",x"c3",x"49",x"73"),
   175 => (x"c0",x"1e",x"71",x"99"),
   176 => (x"87",x"ce",x"fb",x"49"),
   177 => (x"b7",x"c8",x"49",x"73"),
   178 => (x"c1",x"1e",x"71",x"29"),
   179 => (x"87",x"c2",x"fb",x"49"),
   180 => (x"f9",x"c5",x"86",x"c8"),
   181 => (x"e9",x"ed",x"c2",x"87"),
   182 => (x"02",x"9b",x"4b",x"bf"),
   183 => (x"d2",x"c2",x"87",x"dd"),
   184 => (x"c7",x"49",x"bf",x"e4"),
   185 => (x"98",x"70",x"87",x"d6"),
   186 => (x"c0",x"87",x"c4",x"05"),
   187 => (x"c2",x"87",x"d2",x"4b"),
   188 => (x"fb",x"c6",x"49",x"e0"),
   189 => (x"e8",x"d2",x"c2",x"87"),
   190 => (x"c2",x"87",x"c6",x"58"),
   191 => (x"c0",x"48",x"e4",x"d2"),
   192 => (x"c2",x"49",x"73",x"78"),
   193 => (x"87",x"cd",x"05",x"99"),
   194 => (x"e1",x"49",x"eb",x"c3"),
   195 => (x"49",x"70",x"87",x"d6"),
   196 => (x"c2",x"02",x"99",x"c2"),
   197 => (x"73",x"4c",x"fb",x"87"),
   198 => (x"05",x"99",x"c1",x"49"),
   199 => (x"f4",x"c3",x"87",x"cd"),
   200 => (x"87",x"c0",x"e1",x"49"),
   201 => (x"99",x"c2",x"49",x"70"),
   202 => (x"fa",x"87",x"c2",x"02"),
   203 => (x"c8",x"49",x"73",x"4c"),
   204 => (x"87",x"cd",x"05",x"99"),
   205 => (x"e0",x"49",x"f5",x"c3"),
   206 => (x"49",x"70",x"87",x"ea"),
   207 => (x"d4",x"02",x"99",x"c2"),
   208 => (x"f1",x"ed",x"c2",x"87"),
   209 => (x"87",x"c9",x"02",x"bf"),
   210 => (x"c2",x"88",x"c1",x"48"),
   211 => (x"c2",x"58",x"f5",x"ed"),
   212 => (x"c1",x"4c",x"ff",x"87"),
   213 => (x"c4",x"49",x"73",x"4d"),
   214 => (x"87",x"cd",x"05",x"99"),
   215 => (x"e0",x"49",x"f2",x"c3"),
   216 => (x"49",x"70",x"87",x"c2"),
   217 => (x"db",x"02",x"99",x"c2"),
   218 => (x"f1",x"ed",x"c2",x"87"),
   219 => (x"c7",x"48",x"7e",x"bf"),
   220 => (x"cb",x"03",x"a8",x"b7"),
   221 => (x"c1",x"48",x"6e",x"87"),
   222 => (x"f5",x"ed",x"c2",x"80"),
   223 => (x"87",x"c2",x"c0",x"58"),
   224 => (x"4d",x"c1",x"4c",x"fe"),
   225 => (x"ff",x"49",x"fd",x"c3"),
   226 => (x"70",x"87",x"d9",x"df"),
   227 => (x"02",x"99",x"c2",x"49"),
   228 => (x"ed",x"c2",x"87",x"d5"),
   229 => (x"c0",x"02",x"bf",x"f1"),
   230 => (x"ed",x"c2",x"87",x"c9"),
   231 => (x"78",x"c0",x"48",x"f1"),
   232 => (x"fd",x"87",x"c2",x"c0"),
   233 => (x"c3",x"4d",x"c1",x"4c"),
   234 => (x"de",x"ff",x"49",x"fa"),
   235 => (x"49",x"70",x"87",x"f6"),
   236 => (x"d9",x"02",x"99",x"c2"),
   237 => (x"f1",x"ed",x"c2",x"87"),
   238 => (x"b7",x"c7",x"48",x"bf"),
   239 => (x"c9",x"c0",x"03",x"a8"),
   240 => (x"f1",x"ed",x"c2",x"87"),
   241 => (x"c0",x"78",x"c7",x"48"),
   242 => (x"4c",x"fc",x"87",x"c2"),
   243 => (x"b7",x"c0",x"4d",x"c1"),
   244 => (x"d1",x"c0",x"03",x"ac"),
   245 => (x"4a",x"66",x"c4",x"87"),
   246 => (x"6a",x"82",x"d8",x"c1"),
   247 => (x"87",x"c6",x"c0",x"02"),
   248 => (x"49",x"74",x"4b",x"6a"),
   249 => (x"1e",x"c0",x"0f",x"73"),
   250 => (x"c1",x"1e",x"f0",x"c3"),
   251 => (x"dc",x"f7",x"49",x"da"),
   252 => (x"70",x"86",x"c8",x"87"),
   253 => (x"e2",x"c0",x"02",x"98"),
   254 => (x"48",x"a6",x"c8",x"87"),
   255 => (x"bf",x"f1",x"ed",x"c2"),
   256 => (x"49",x"66",x"c8",x"78"),
   257 => (x"66",x"c4",x"91",x"cb"),
   258 => (x"70",x"80",x"71",x"48"),
   259 => (x"02",x"bf",x"6e",x"7e"),
   260 => (x"6e",x"87",x"c8",x"c0"),
   261 => (x"66",x"c8",x"4b",x"bf"),
   262 => (x"75",x"0f",x"73",x"49"),
   263 => (x"c8",x"c0",x"02",x"9d"),
   264 => (x"f1",x"ed",x"c2",x"87"),
   265 => (x"ca",x"f3",x"49",x"bf"),
   266 => (x"ec",x"d2",x"c2",x"87"),
   267 => (x"dd",x"c0",x"02",x"bf"),
   268 => (x"c7",x"c2",x"49",x"87"),
   269 => (x"02",x"98",x"70",x"87"),
   270 => (x"c2",x"87",x"d3",x"c0"),
   271 => (x"49",x"bf",x"f1",x"ed"),
   272 => (x"c0",x"87",x"f0",x"f2"),
   273 => (x"87",x"d0",x"f4",x"49"),
   274 => (x"48",x"ec",x"d2",x"c2"),
   275 => (x"8e",x"f4",x"78",x"c0"),
   276 => (x"0e",x"87",x"ea",x"f3"),
   277 => (x"5d",x"5c",x"5b",x"5e"),
   278 => (x"4c",x"71",x"1e",x"0e"),
   279 => (x"bf",x"ed",x"ed",x"c2"),
   280 => (x"a1",x"cd",x"c1",x"49"),
   281 => (x"81",x"d1",x"c1",x"4d"),
   282 => (x"9c",x"74",x"7e",x"69"),
   283 => (x"c4",x"87",x"cf",x"02"),
   284 => (x"7b",x"74",x"4b",x"a5"),
   285 => (x"bf",x"ed",x"ed",x"c2"),
   286 => (x"87",x"c9",x"f3",x"49"),
   287 => (x"9c",x"74",x"7b",x"6e"),
   288 => (x"c0",x"87",x"c4",x"05"),
   289 => (x"c1",x"87",x"c2",x"4b"),
   290 => (x"f3",x"49",x"73",x"4b"),
   291 => (x"66",x"d4",x"87",x"ca"),
   292 => (x"49",x"87",x"c7",x"02"),
   293 => (x"4a",x"70",x"87",x"da"),
   294 => (x"4a",x"c0",x"87",x"c2"),
   295 => (x"5a",x"f0",x"d2",x"c2"),
   296 => (x"87",x"d9",x"f2",x"26"),
   297 => (x"00",x"00",x"00",x"00"),
   298 => (x"00",x"00",x"00",x"00"),
   299 => (x"00",x"00",x"00",x"00"),
   300 => (x"ff",x"4a",x"71",x"1e"),
   301 => (x"72",x"49",x"bf",x"c8"),
   302 => (x"4f",x"26",x"48",x"a1"),
   303 => (x"bf",x"c8",x"ff",x"1e"),
   304 => (x"c0",x"c0",x"fe",x"89"),
   305 => (x"a9",x"c0",x"c0",x"c0"),
   306 => (x"c0",x"87",x"c4",x"01"),
   307 => (x"c1",x"87",x"c2",x"4a"),
   308 => (x"26",x"48",x"72",x"4a"),
   309 => (x"5b",x"5e",x"0e",x"4f"),
   310 => (x"71",x"0e",x"5d",x"5c"),
   311 => (x"4c",x"d4",x"ff",x"4b"),
   312 => (x"c0",x"48",x"66",x"d0"),
   313 => (x"ff",x"49",x"d6",x"78"),
   314 => (x"c3",x"87",x"f1",x"db"),
   315 => (x"49",x"6c",x"7c",x"ff"),
   316 => (x"71",x"99",x"ff",x"c3"),
   317 => (x"f0",x"c3",x"49",x"4d"),
   318 => (x"a9",x"e0",x"c1",x"99"),
   319 => (x"c3",x"87",x"cb",x"05"),
   320 => (x"48",x"6c",x"7c",x"ff"),
   321 => (x"66",x"d0",x"98",x"c3"),
   322 => (x"ff",x"c3",x"78",x"08"),
   323 => (x"49",x"4a",x"6c",x"7c"),
   324 => (x"ff",x"c3",x"31",x"c8"),
   325 => (x"71",x"4a",x"6c",x"7c"),
   326 => (x"c8",x"49",x"72",x"b2"),
   327 => (x"7c",x"ff",x"c3",x"31"),
   328 => (x"b2",x"71",x"4a",x"6c"),
   329 => (x"31",x"c8",x"49",x"72"),
   330 => (x"6c",x"7c",x"ff",x"c3"),
   331 => (x"ff",x"b2",x"71",x"4a"),
   332 => (x"e0",x"c0",x"48",x"d0"),
   333 => (x"02",x"9b",x"73",x"78"),
   334 => (x"7b",x"72",x"87",x"c2"),
   335 => (x"4d",x"26",x"48",x"75"),
   336 => (x"4b",x"26",x"4c",x"26"),
   337 => (x"26",x"1e",x"4f",x"26"),
   338 => (x"5b",x"5e",x"0e",x"4f"),
   339 => (x"86",x"f8",x"0e",x"5c"),
   340 => (x"a6",x"c8",x"1e",x"76"),
   341 => (x"87",x"fd",x"fd",x"49"),
   342 => (x"4b",x"70",x"86",x"c4"),
   343 => (x"a8",x"c2",x"48",x"6e"),
   344 => (x"87",x"f0",x"c2",x"03"),
   345 => (x"f0",x"c3",x"4a",x"73"),
   346 => (x"aa",x"d0",x"c1",x"9a"),
   347 => (x"c1",x"87",x"c7",x"02"),
   348 => (x"c2",x"05",x"aa",x"e0"),
   349 => (x"49",x"73",x"87",x"de"),
   350 => (x"c3",x"02",x"99",x"c8"),
   351 => (x"87",x"c6",x"ff",x"87"),
   352 => (x"9c",x"c3",x"4c",x"73"),
   353 => (x"c1",x"05",x"ac",x"c2"),
   354 => (x"66",x"c4",x"87",x"c2"),
   355 => (x"71",x"31",x"c9",x"49"),
   356 => (x"4a",x"66",x"c4",x"1e"),
   357 => (x"ed",x"c2",x"92",x"d4"),
   358 => (x"81",x"72",x"49",x"f5"),
   359 => (x"87",x"c0",x"d1",x"fe"),
   360 => (x"d8",x"ff",x"49",x"d8"),
   361 => (x"c0",x"c8",x"87",x"f6"),
   362 => (x"d2",x"dc",x"c2",x"1e"),
   363 => (x"fb",x"ec",x"fd",x"49"),
   364 => (x"48",x"d0",x"ff",x"87"),
   365 => (x"c2",x"78",x"e0",x"c0"),
   366 => (x"cc",x"1e",x"d2",x"dc"),
   367 => (x"92",x"d4",x"4a",x"66"),
   368 => (x"49",x"f5",x"ed",x"c2"),
   369 => (x"cf",x"fe",x"81",x"72"),
   370 => (x"86",x"cc",x"87",x"c7"),
   371 => (x"c1",x"05",x"ac",x"c1"),
   372 => (x"66",x"c4",x"87",x"c2"),
   373 => (x"71",x"31",x"c9",x"49"),
   374 => (x"4a",x"66",x"c4",x"1e"),
   375 => (x"ed",x"c2",x"92",x"d4"),
   376 => (x"81",x"72",x"49",x"f5"),
   377 => (x"87",x"f8",x"cf",x"fe"),
   378 => (x"1e",x"d2",x"dc",x"c2"),
   379 => (x"d4",x"4a",x"66",x"c8"),
   380 => (x"f5",x"ed",x"c2",x"92"),
   381 => (x"fe",x"81",x"72",x"49"),
   382 => (x"d7",x"87",x"c7",x"cd"),
   383 => (x"db",x"d7",x"ff",x"49"),
   384 => (x"1e",x"c0",x"c8",x"87"),
   385 => (x"49",x"d2",x"dc",x"c2"),
   386 => (x"87",x"f9",x"ea",x"fd"),
   387 => (x"d0",x"ff",x"86",x"cc"),
   388 => (x"78",x"e0",x"c0",x"48"),
   389 => (x"e7",x"fc",x"8e",x"f8"),
   390 => (x"5b",x"5e",x"0e",x"87"),
   391 => (x"1e",x"0e",x"5d",x"5c"),
   392 => (x"d4",x"ff",x"4d",x"71"),
   393 => (x"7e",x"66",x"d4",x"4c"),
   394 => (x"a8",x"b7",x"c3",x"48"),
   395 => (x"c0",x"87",x"c5",x"06"),
   396 => (x"87",x"e2",x"c1",x"48"),
   397 => (x"dd",x"fe",x"49",x"75"),
   398 => (x"1e",x"75",x"87",x"fb"),
   399 => (x"d4",x"4b",x"66",x"c4"),
   400 => (x"f5",x"ed",x"c2",x"93"),
   401 => (x"fe",x"49",x"73",x"83"),
   402 => (x"c8",x"87",x"e2",x"c8"),
   403 => (x"ff",x"4b",x"6b",x"83"),
   404 => (x"e1",x"c8",x"48",x"d0"),
   405 => (x"73",x"7c",x"dd",x"78"),
   406 => (x"99",x"ff",x"c3",x"49"),
   407 => (x"49",x"73",x"7c",x"71"),
   408 => (x"c3",x"29",x"b7",x"c8"),
   409 => (x"7c",x"71",x"99",x"ff"),
   410 => (x"b7",x"d0",x"49",x"73"),
   411 => (x"99",x"ff",x"c3",x"29"),
   412 => (x"49",x"73",x"7c",x"71"),
   413 => (x"71",x"29",x"b7",x"d8"),
   414 => (x"7c",x"7c",x"c0",x"7c"),
   415 => (x"7c",x"7c",x"7c",x"7c"),
   416 => (x"7c",x"7c",x"7c",x"7c"),
   417 => (x"e0",x"c0",x"7c",x"7c"),
   418 => (x"1e",x"66",x"c4",x"78"),
   419 => (x"d5",x"ff",x"49",x"dc"),
   420 => (x"86",x"c8",x"87",x"ef"),
   421 => (x"fa",x"26",x"48",x"73"),
   422 => (x"c2",x"1e",x"87",x"e4"),
   423 => (x"49",x"bf",x"e8",x"db"),
   424 => (x"db",x"c2",x"b9",x"c1"),
   425 => (x"d4",x"ff",x"59",x"ec"),
   426 => (x"78",x"ff",x"c3",x"48"),
   427 => (x"c8",x"48",x"d0",x"ff"),
   428 => (x"d4",x"ff",x"78",x"e1"),
   429 => (x"c4",x"78",x"c1",x"48"),
   430 => (x"ff",x"78",x"71",x"31"),
   431 => (x"e0",x"c0",x"48",x"d0"),
   432 => (x"1e",x"4f",x"26",x"78"),
   433 => (x"1e",x"dc",x"db",x"c2"),
   434 => (x"49",x"c8",x"e9",x"c2"),
   435 => (x"87",x"dd",x"c6",x"fe"),
   436 => (x"98",x"70",x"86",x"c4"),
   437 => (x"ff",x"87",x"c3",x"02"),
   438 => (x"4f",x"26",x"87",x"c0"),
   439 => (x"48",x"4b",x"35",x"31"),
   440 => (x"20",x"20",x"20",x"5a"),
   441 => (x"00",x"47",x"46",x"43"),
   442 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

