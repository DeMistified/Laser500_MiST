library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"e0eec287",
    12 => x"86c0c64e",
    13 => x"49e0eec2",
    14 => x"48ecdbc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087f0e1",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"4a711e4f",
    50 => x"484966c4",
    51 => x"a6c888c1",
    52 => x"02997158",
    53 => x"481287d4",
    54 => x"7808d4ff",
    55 => x"484966c4",
    56 => x"a6c888c1",
    57 => x"05997158",
    58 => x"4f2687ec",
    59 => x"c44a711e",
    60 => x"c1484966",
    61 => x"58a6c888",
    62 => x"d6029971",
    63 => x"48d4ff87",
    64 => x"6878ffc3",
    65 => x"4966c452",
    66 => x"c888c148",
    67 => x"997158a6",
    68 => x"2687ea05",
    69 => x"1e731e4f",
    70 => x"c34bd4ff",
    71 => x"4a6b7bff",
    72 => x"6b7bffc3",
    73 => x"7232c849",
    74 => x"7bffc3b1",
    75 => x"31c84a6b",
    76 => x"ffc3b271",
    77 => x"c8496b7b",
    78 => x"71b17232",
    79 => x"2687c448",
    80 => x"264c264d",
    81 => x"0e4f264b",
    82 => x"5d5c5b5e",
    83 => x"ff4a710e",
    84 => x"49724cd4",
    85 => x"7199ffc3",
    86 => x"ecdbc27c",
    87 => x"87c805bf",
    88 => x"c94866d0",
    89 => x"58a6d430",
    90 => x"d84966d0",
    91 => x"99ffc329",
    92 => x"66d07c71",
    93 => x"c329d049",
    94 => x"7c7199ff",
    95 => x"c84966d0",
    96 => x"99ffc329",
    97 => x"66d07c71",
    98 => x"99ffc349",
    99 => x"49727c71",
   100 => x"ffc329d0",
   101 => x"6c7c7199",
   102 => x"fff0c94b",
   103 => x"abffc34d",
   104 => x"c387d005",
   105 => x"4b6c7cff",
   106 => x"c6028dc1",
   107 => x"abffc387",
   108 => x"7387f002",
   109 => x"87c7fe48",
   110 => x"ff49c01e",
   111 => x"ffc348d4",
   112 => x"c381c178",
   113 => x"04a9b7c8",
   114 => x"4f2687f1",
   115 => x"e71e731e",
   116 => x"dff8c487",
   117 => x"c01ec04b",
   118 => x"f7c1f0ff",
   119 => x"87e7fd49",
   120 => x"a8c186c4",
   121 => x"87eac005",
   122 => x"c348d4ff",
   123 => x"c0c178ff",
   124 => x"c0c0c0c0",
   125 => x"f0e1c01e",
   126 => x"fd49e9c1",
   127 => x"86c487c9",
   128 => x"ca059870",
   129 => x"48d4ff87",
   130 => x"c178ffc3",
   131 => x"fe87cb48",
   132 => x"8bc187e6",
   133 => x"87fdfe05",
   134 => x"e6fc48c0",
   135 => x"1e731e87",
   136 => x"c348d4ff",
   137 => x"4bd378ff",
   138 => x"ffc01ec0",
   139 => x"49c1c1f0",
   140 => x"c487d4fc",
   141 => x"05987086",
   142 => x"d4ff87ca",
   143 => x"78ffc348",
   144 => x"87cb48c1",
   145 => x"c187f1fd",
   146 => x"dbff058b",
   147 => x"fb48c087",
   148 => x"5e0e87f1",
   149 => x"ff0e5c5b",
   150 => x"dbfd4cd4",
   151 => x"1eeac687",
   152 => x"c1f0e1c0",
   153 => x"defb49c8",
   154 => x"c186c487",
   155 => x"87c802a8",
   156 => x"c087eafe",
   157 => x"87e2c148",
   158 => x"7087dafa",
   159 => x"ffffcf49",
   160 => x"a9eac699",
   161 => x"fe87c802",
   162 => x"48c087d3",
   163 => x"c387cbc1",
   164 => x"f1c07cff",
   165 => x"87f4fc4b",
   166 => x"c0029870",
   167 => x"1ec087eb",
   168 => x"c1f0ffc0",
   169 => x"defa49fa",
   170 => x"7086c487",
   171 => x"87d90598",
   172 => x"6c7cffc3",
   173 => x"7cffc349",
   174 => x"c17c7c7c",
   175 => x"c40299c0",
   176 => x"d548c187",
   177 => x"d148c087",
   178 => x"05abc287",
   179 => x"48c087c4",
   180 => x"8bc187c8",
   181 => x"87fdfe05",
   182 => x"e4f948c0",
   183 => x"1e731e87",
   184 => x"48ecdbc2",
   185 => x"4bc778c1",
   186 => x"c248d0ff",
   187 => x"87c8fb78",
   188 => x"c348d0ff",
   189 => x"c01ec078",
   190 => x"c0c1d0e5",
   191 => x"87c7f949",
   192 => x"a8c186c4",
   193 => x"4b87c105",
   194 => x"c505abc2",
   195 => x"c048c087",
   196 => x"8bc187f9",
   197 => x"87d0ff05",
   198 => x"c287f7fc",
   199 => x"7058f0db",
   200 => x"87cd0598",
   201 => x"ffc01ec1",
   202 => x"49d0c1f0",
   203 => x"c487d8f8",
   204 => x"48d4ff86",
   205 => x"c478ffc3",
   206 => x"dbc287de",
   207 => x"d0ff58f4",
   208 => x"ff78c248",
   209 => x"ffc348d4",
   210 => x"f748c178",
   211 => x"5e0e87f5",
   212 => x"0e5d5c5b",
   213 => x"ffc34a71",
   214 => x"4cd4ff4d",
   215 => x"d0ff7c75",
   216 => x"78c3c448",
   217 => x"1e727c75",
   218 => x"c1f0ffc0",
   219 => x"d6f749d8",
   220 => x"7086c487",
   221 => x"87c50298",
   222 => x"f0c048c1",
   223 => x"c37c7587",
   224 => x"c0c87cfe",
   225 => x"4966d41e",
   226 => x"c487faf4",
   227 => x"757c7586",
   228 => x"d87c757c",
   229 => x"754be0da",
   230 => x"99496c7c",
   231 => x"c187c505",
   232 => x"87f3058b",
   233 => x"d0ff7c75",
   234 => x"c078c248",
   235 => x"87cff648",
   236 => x"5c5b5e0e",
   237 => x"4b710e5d",
   238 => x"eec54cc0",
   239 => x"ff4adfcd",
   240 => x"ffc348d4",
   241 => x"c3496878",
   242 => x"c005a9fe",
   243 => x"4d7087fd",
   244 => x"cc029b73",
   245 => x"1e66d087",
   246 => x"cff44973",
   247 => x"d686c487",
   248 => x"48d0ff87",
   249 => x"c378d1c4",
   250 => x"66d07dff",
   251 => x"d488c148",
   252 => x"987058a6",
   253 => x"ff87f005",
   254 => x"ffc348d4",
   255 => x"9b737878",
   256 => x"ff87c505",
   257 => x"78d048d0",
   258 => x"c14c4ac1",
   259 => x"eefe058a",
   260 => x"f4487487",
   261 => x"731e87e9",
   262 => x"c04a711e",
   263 => x"48d4ff4b",
   264 => x"ff78ffc3",
   265 => x"c3c448d0",
   266 => x"48d4ff78",
   267 => x"7278ffc3",
   268 => x"f0ffc01e",
   269 => x"f449d1c1",
   270 => x"86c487cd",
   271 => x"d2059870",
   272 => x"1ec0c887",
   273 => x"fd4966cc",
   274 => x"86c487e6",
   275 => x"d0ff4b70",
   276 => x"7378c248",
   277 => x"87ebf348",
   278 => x"5c5b5e0e",
   279 => x"1ec00e5d",
   280 => x"c1f0ffc0",
   281 => x"def349c9",
   282 => x"c21ed287",
   283 => x"fc49f4db",
   284 => x"86c887fe",
   285 => x"84c14cc0",
   286 => x"04acb7d2",
   287 => x"dbc287f8",
   288 => x"49bf97f4",
   289 => x"c199c0c3",
   290 => x"c005a9c0",
   291 => x"dbc287e7",
   292 => x"49bf97fb",
   293 => x"dbc231d0",
   294 => x"4abf97fc",
   295 => x"b17232c8",
   296 => x"97fddbc2",
   297 => x"71b14abf",
   298 => x"ffffcf4c",
   299 => x"84c19cff",
   300 => x"e7c134ca",
   301 => x"fddbc287",
   302 => x"c149bf97",
   303 => x"c299c631",
   304 => x"bf97fedb",
   305 => x"2ab7c74a",
   306 => x"dbc2b172",
   307 => x"4abf97f9",
   308 => x"c29dcf4d",
   309 => x"bf97fadb",
   310 => x"ca9ac34a",
   311 => x"fbdbc232",
   312 => x"c24bbf97",
   313 => x"c2b27333",
   314 => x"bf97fcdb",
   315 => x"9bc0c34b",
   316 => x"732bb7c6",
   317 => x"c181c2b2",
   318 => x"70307148",
   319 => x"7548c149",
   320 => x"724d7030",
   321 => x"7184c14c",
   322 => x"b7c0c894",
   323 => x"87cc06ad",
   324 => x"2db734c1",
   325 => x"adb7c0c8",
   326 => x"87f4ff01",
   327 => x"def04874",
   328 => x"5b5e0e87",
   329 => x"f80e5d5c",
   330 => x"dae4c286",
   331 => x"c278c048",
   332 => x"c01ed2dc",
   333 => x"87defb49",
   334 => x"987086c4",
   335 => x"c087c505",
   336 => x"87cec948",
   337 => x"7ec14dc0",
   338 => x"bfc0f3c0",
   339 => x"c8ddc249",
   340 => x"4bc8714a",
   341 => x"7087d3ec",
   342 => x"87c20598",
   343 => x"f2c07ec0",
   344 => x"c249bffc",
   345 => x"714ae4dd",
   346 => x"fdeb4bc8",
   347 => x"05987087",
   348 => x"7ec087c2",
   349 => x"fdc0026e",
   350 => x"d8e3c287",
   351 => x"e4c24dbf",
   352 => x"7ebf9fd0",
   353 => x"ead6c548",
   354 => x"87c705a8",
   355 => x"bfd8e3c2",
   356 => x"6e87ce4d",
   357 => x"d5e9ca48",
   358 => x"87c502a8",
   359 => x"f1c748c0",
   360 => x"d2dcc287",
   361 => x"f949751e",
   362 => x"86c487ec",
   363 => x"c5059870",
   364 => x"c748c087",
   365 => x"f2c087dc",
   366 => x"c249bffc",
   367 => x"714ae4dd",
   368 => x"e5ea4bc8",
   369 => x"05987087",
   370 => x"e4c287c8",
   371 => x"78c148da",
   372 => x"f3c087da",
   373 => x"c249bfc0",
   374 => x"714ac8dd",
   375 => x"c9ea4bc8",
   376 => x"02987087",
   377 => x"c087c5c0",
   378 => x"87e6c648",
   379 => x"97d0e4c2",
   380 => x"d5c149bf",
   381 => x"cdc005a9",
   382 => x"d1e4c287",
   383 => x"c249bf97",
   384 => x"c002a9ea",
   385 => x"48c087c5",
   386 => x"c287c7c6",
   387 => x"bf97d2dc",
   388 => x"e9c3487e",
   389 => x"cec002a8",
   390 => x"c3486e87",
   391 => x"c002a8eb",
   392 => x"48c087c5",
   393 => x"c287ebc5",
   394 => x"bf97dddc",
   395 => x"c0059949",
   396 => x"dcc287cc",
   397 => x"49bf97de",
   398 => x"c002a9c2",
   399 => x"48c087c5",
   400 => x"c287cfc5",
   401 => x"bf97dfdc",
   402 => x"d6e4c248",
   403 => x"484c7058",
   404 => x"e4c288c1",
   405 => x"dcc258da",
   406 => x"49bf97e0",
   407 => x"dcc28175",
   408 => x"4abf97e1",
   409 => x"a17232c8",
   410 => x"e7e8c27e",
   411 => x"c2786e48",
   412 => x"bf97e2dc",
   413 => x"58a6c848",
   414 => x"bfdae4c2",
   415 => x"87d4c202",
   416 => x"bffcf2c0",
   417 => x"e4ddc249",
   418 => x"4bc8714a",
   419 => x"7087dbe7",
   420 => x"c5c00298",
   421 => x"c348c087",
   422 => x"e4c287f8",
   423 => x"c24cbfd2",
   424 => x"c25cfbe8",
   425 => x"bf97f7dc",
   426 => x"c231c849",
   427 => x"bf97f6dc",
   428 => x"c249a14a",
   429 => x"bf97f8dc",
   430 => x"7232d04a",
   431 => x"dcc249a1",
   432 => x"4abf97f9",
   433 => x"a17232d8",
   434 => x"9166c449",
   435 => x"bfe7e8c2",
   436 => x"efe8c281",
   437 => x"ffdcc259",
   438 => x"c84abf97",
   439 => x"fedcc232",
   440 => x"a24bbf97",
   441 => x"c0ddc24a",
   442 => x"d04bbf97",
   443 => x"4aa27333",
   444 => x"97c1ddc2",
   445 => x"9bcf4bbf",
   446 => x"a27333d8",
   447 => x"f3e8c24a",
   448 => x"efe8c25a",
   449 => x"8ac24abf",
   450 => x"e8c29274",
   451 => x"a17248f3",
   452 => x"87cac178",
   453 => x"97e4dcc2",
   454 => x"31c849bf",
   455 => x"97e3dcc2",
   456 => x"49a14abf",
   457 => x"59e2e4c2",
   458 => x"bfdee4c2",
   459 => x"c731c549",
   460 => x"29c981ff",
   461 => x"59fbe8c2",
   462 => x"97e9dcc2",
   463 => x"32c84abf",
   464 => x"97e8dcc2",
   465 => x"4aa24bbf",
   466 => x"6e9266c4",
   467 => x"f7e8c282",
   468 => x"efe8c25a",
   469 => x"c278c048",
   470 => x"7248ebe8",
   471 => x"e8c278a1",
   472 => x"e8c248fb",
   473 => x"c278bfef",
   474 => x"c248ffe8",
   475 => x"78bff3e8",
   476 => x"bfdae4c2",
   477 => x"87c9c002",
   478 => x"30c44874",
   479 => x"c9c07e70",
   480 => x"f7e8c287",
   481 => x"30c448bf",
   482 => x"e4c27e70",
   483 => x"786e48de",
   484 => x"8ef848c1",
   485 => x"4c264d26",
   486 => x"4f264b26",
   487 => x"5c5b5e0e",
   488 => x"4a710e5d",
   489 => x"bfdae4c2",
   490 => x"7287cb02",
   491 => x"722bc74b",
   492 => x"9cffc14c",
   493 => x"4b7287c9",
   494 => x"4c722bc8",
   495 => x"c29cffc3",
   496 => x"83bfe7e8",
   497 => x"bff8f2c0",
   498 => x"87d902ab",
   499 => x"5bfcf2c0",
   500 => x"1ed2dcc2",
   501 => x"fdf04973",
   502 => x"7086c487",
   503 => x"87c50598",
   504 => x"e6c048c0",
   505 => x"dae4c287",
   506 => x"87d202bf",
   507 => x"91c44974",
   508 => x"81d2dcc2",
   509 => x"ffcf4d69",
   510 => x"9dffffff",
   511 => x"497487cb",
   512 => x"dcc291c2",
   513 => x"699f81d2",
   514 => x"fe48754d",
   515 => x"5e0e87c6",
   516 => x"0e5d5c5b",
   517 => x"c04d711e",
   518 => x"ca49c11e",
   519 => x"86c487ff",
   520 => x"029c4c70",
   521 => x"c287c0c1",
   522 => x"754ae2e4",
   523 => x"87dfe049",
   524 => x"c0029870",
   525 => x"4a7487f1",
   526 => x"4bcb4975",
   527 => x"7087c5e1",
   528 => x"e2c00298",
   529 => x"741ec087",
   530 => x"87c7029c",
   531 => x"c048a6c4",
   532 => x"c487c578",
   533 => x"78c148a6",
   534 => x"c94966c4",
   535 => x"86c487ff",
   536 => x"059c4c70",
   537 => x"7487c0ff",
   538 => x"e7fc2648",
   539 => x"5b5e0e87",
   540 => x"1e0e5d5c",
   541 => x"059b4b71",
   542 => x"48c087c5",
   543 => x"c887e5c1",
   544 => x"7dc04da3",
   545 => x"c70266d4",
   546 => x"9766d487",
   547 => x"87c505bf",
   548 => x"cfc148c0",
   549 => x"4966d487",
   550 => x"7087f3fd",
   551 => x"c1029c4c",
   552 => x"a4dc87c0",
   553 => x"da7d6949",
   554 => x"a3c449a4",
   555 => x"7a699f4a",
   556 => x"bfdae4c2",
   557 => x"d487d202",
   558 => x"699f49a4",
   559 => x"ffffc049",
   560 => x"d0487199",
   561 => x"c27e7030",
   562 => x"6e7ec087",
   563 => x"806a4849",
   564 => x"7bc07a70",
   565 => x"6a49a3cc",
   566 => x"49a3d079",
   567 => x"48c179c0",
   568 => x"48c087c2",
   569 => x"87ecfa26",
   570 => x"5c5b5e0e",
   571 => x"4c710e5d",
   572 => x"cac1029c",
   573 => x"49a4c887",
   574 => x"c2c10269",
   575 => x"4a66d087",
   576 => x"d482496c",
   577 => x"66d05aa6",
   578 => x"e4c2b94d",
   579 => x"ff4abfd6",
   580 => x"719972ba",
   581 => x"e4c00299",
   582 => x"4ba4c487",
   583 => x"fbf9496b",
   584 => x"c27b7087",
   585 => x"49bfd2e4",
   586 => x"7c71816c",
   587 => x"e4c2b975",
   588 => x"ff4abfd6",
   589 => x"719972ba",
   590 => x"dcff0599",
   591 => x"f97c7587",
   592 => x"731e87d2",
   593 => x"9b4b711e",
   594 => x"c887c702",
   595 => x"056949a3",
   596 => x"48c087c5",
   597 => x"c287f7c0",
   598 => x"4abfebe8",
   599 => x"6949a3c4",
   600 => x"c289c249",
   601 => x"91bfd2e4",
   602 => x"c24aa271",
   603 => x"49bfd6e4",
   604 => x"a271996b",
   605 => x"fcf2c04a",
   606 => x"1e66c85a",
   607 => x"d5ea4972",
   608 => x"7086c487",
   609 => x"87c40598",
   610 => x"87c248c0",
   611 => x"c7f848c1",
   612 => x"1e731e87",
   613 => x"029b4b71",
   614 => x"a3c887c7",
   615 => x"c5056949",
   616 => x"c048c087",
   617 => x"e8c287f7",
   618 => x"c44abfeb",
   619 => x"496949a3",
   620 => x"e4c289c2",
   621 => x"7191bfd2",
   622 => x"e4c24aa2",
   623 => x"6b49bfd6",
   624 => x"4aa27199",
   625 => x"5afcf2c0",
   626 => x"721e66c8",
   627 => x"87fee549",
   628 => x"987086c4",
   629 => x"c087c405",
   630 => x"c187c248",
   631 => x"87f8f648",
   632 => x"5c5b5e0e",
   633 => x"711e0e5d",
   634 => x"4c66d44b",
   635 => x"9b732cc9",
   636 => x"87cfc102",
   637 => x"6949a3c8",
   638 => x"87c7c102",
   639 => x"d44da3d0",
   640 => x"e4c27d66",
   641 => x"ff49bfd6",
   642 => x"994a6bb9",
   643 => x"03ac717e",
   644 => x"7bc087cd",
   645 => x"4aa3cc7d",
   646 => x"6a49a3c4",
   647 => x"7287c279",
   648 => x"029c748c",
   649 => x"1e4987dd",
   650 => x"fbfa4973",
   651 => x"d486c487",
   652 => x"ffc74966",
   653 => x"87cb0299",
   654 => x"1ed2dcc2",
   655 => x"c1fc4973",
   656 => x"2686c487",
   657 => x"1e87cdf5",
   658 => x"4b711e73",
   659 => x"e4c0029b",
   660 => x"ffe8c287",
   661 => x"c24a735b",
   662 => x"d2e4c28a",
   663 => x"c29249bf",
   664 => x"48bfebe8",
   665 => x"e9c28072",
   666 => x"487158c3",
   667 => x"e4c230c4",
   668 => x"edc058e2",
   669 => x"fbe8c287",
   670 => x"efe8c248",
   671 => x"e8c278bf",
   672 => x"e8c248ff",
   673 => x"c278bff3",
   674 => x"02bfdae4",
   675 => x"e4c287c9",
   676 => x"c449bfd2",
   677 => x"c287c731",
   678 => x"49bff7e8",
   679 => x"e4c231c4",
   680 => x"f3f359e2",
   681 => x"5b5e0e87",
   682 => x"4a710e5c",
   683 => x"9a724bc0",
   684 => x"87e1c002",
   685 => x"9f49a2da",
   686 => x"e4c24b69",
   687 => x"cf02bfda",
   688 => x"49a2d487",
   689 => x"4c49699f",
   690 => x"9cffffc0",
   691 => x"87c234d0",
   692 => x"49744cc0",
   693 => x"fd4973b3",
   694 => x"f9f287ed",
   695 => x"5b5e0e87",
   696 => x"f40e5d5c",
   697 => x"c04a7186",
   698 => x"029a727e",
   699 => x"dcc287d8",
   700 => x"78c048ce",
   701 => x"48c6dcc2",
   702 => x"bfffe8c2",
   703 => x"cadcc278",
   704 => x"fbe8c248",
   705 => x"e4c278bf",
   706 => x"50c048ef",
   707 => x"bfdee4c2",
   708 => x"cedcc249",
   709 => x"aa714abf",
   710 => x"87c9c403",
   711 => x"99cf4972",
   712 => x"87e9c005",
   713 => x"48f8f2c0",
   714 => x"bfc6dcc2",
   715 => x"d2dcc278",
   716 => x"c6dcc21e",
   717 => x"dcc249bf",
   718 => x"a1c148c6",
   719 => x"d5e37178",
   720 => x"c086c487",
   721 => x"c248f4f2",
   722 => x"cc78d2dc",
   723 => x"f4f2c087",
   724 => x"e0c048bf",
   725 => x"f8f2c080",
   726 => x"cedcc258",
   727 => x"80c148bf",
   728 => x"58d2dcc2",
   729 => x"000cb427",
   730 => x"bf97bf00",
   731 => x"c2029d4d",
   732 => x"e5c387e3",
   733 => x"dcc202ad",
   734 => x"f4f2c087",
   735 => x"a3cb4bbf",
   736 => x"cf4c1149",
   737 => x"d2c105ac",
   738 => x"df497587",
   739 => x"cd89c199",
   740 => x"e2e4c291",
   741 => x"4aa3c181",
   742 => x"a3c35112",
   743 => x"c551124a",
   744 => x"51124aa3",
   745 => x"124aa3c7",
   746 => x"4aa3c951",
   747 => x"a3ce5112",
   748 => x"d051124a",
   749 => x"51124aa3",
   750 => x"124aa3d2",
   751 => x"4aa3d451",
   752 => x"a3d65112",
   753 => x"d851124a",
   754 => x"51124aa3",
   755 => x"124aa3dc",
   756 => x"4aa3de51",
   757 => x"7ec15112",
   758 => x"7487fac0",
   759 => x"0599c849",
   760 => x"7487ebc0",
   761 => x"0599d049",
   762 => x"66dc87d1",
   763 => x"87cbc002",
   764 => x"66dc4973",
   765 => x"0298700f",
   766 => x"6e87d3c0",
   767 => x"87c6c005",
   768 => x"48e2e4c2",
   769 => x"f2c050c0",
   770 => x"c248bff4",
   771 => x"e4c287e1",
   772 => x"50c048ef",
   773 => x"dee4c27e",
   774 => x"dcc249bf",
   775 => x"714abfce",
   776 => x"f7fb04aa",
   777 => x"ffe8c287",
   778 => x"c8c005bf",
   779 => x"dae4c287",
   780 => x"f8c102bf",
   781 => x"cadcc287",
   782 => x"dfed49bf",
   783 => x"c2497087",
   784 => x"c459cedc",
   785 => x"dcc248a6",
   786 => x"c278bfca",
   787 => x"02bfdae4",
   788 => x"c487d8c0",
   789 => x"ffcf4966",
   790 => x"99f8ffff",
   791 => x"c5c002a9",
   792 => x"c04cc087",
   793 => x"4cc187e1",
   794 => x"c487dcc0",
   795 => x"ffcf4966",
   796 => x"02a999f8",
   797 => x"c887c8c0",
   798 => x"78c048a6",
   799 => x"c887c5c0",
   800 => x"78c148a6",
   801 => x"744c66c8",
   802 => x"e0c0059c",
   803 => x"4966c487",
   804 => x"e4c289c2",
   805 => x"914abfd2",
   806 => x"bfebe8c2",
   807 => x"c6dcc24a",
   808 => x"78a17248",
   809 => x"48cedcc2",
   810 => x"dff978c0",
   811 => x"f448c087",
   812 => x"87e0eb8e",
   813 => x"00000000",
   814 => x"ffffffff",
   815 => x"00000cc4",
   816 => x"00000ccd",
   817 => x"33544146",
   818 => x"20202032",
   819 => x"54414600",
   820 => x"20203631",
   821 => x"ff1e0020",
   822 => x"ffc348d4",
   823 => x"26486878",
   824 => x"d4ff1e4f",
   825 => x"78ffc348",
   826 => x"c848d0ff",
   827 => x"d4ff78e1",
   828 => x"c278d448",
   829 => x"ff48c3e9",
   830 => x"2650bfd4",
   831 => x"d0ff1e4f",
   832 => x"78e0c048",
   833 => x"ff1e4f26",
   834 => x"497087cc",
   835 => x"87c60299",
   836 => x"05a9fbc0",
   837 => x"487187f1",
   838 => x"5e0e4f26",
   839 => x"710e5c5b",
   840 => x"fe4cc04b",
   841 => x"497087f0",
   842 => x"f9c00299",
   843 => x"a9ecc087",
   844 => x"87f2c002",
   845 => x"02a9fbc0",
   846 => x"cc87ebc0",
   847 => x"03acb766",
   848 => x"66d087c7",
   849 => x"7187c202",
   850 => x"02997153",
   851 => x"84c187c2",
   852 => x"7087c3fe",
   853 => x"cd029949",
   854 => x"a9ecc087",
   855 => x"c087c702",
   856 => x"ff05a9fb",
   857 => x"66d087d5",
   858 => x"c087c302",
   859 => x"ecc07b97",
   860 => x"87c405a9",
   861 => x"87c54a74",
   862 => x"0ac04a74",
   863 => x"c248728a",
   864 => x"264d2687",
   865 => x"264b264c",
   866 => x"c9fd1e4f",
   867 => x"c0497087",
   868 => x"04a9b7f0",
   869 => x"f9c087ca",
   870 => x"c301a9b7",
   871 => x"89f0c087",
   872 => x"a9b7c1c1",
   873 => x"c187ca04",
   874 => x"01a9b7da",
   875 => x"f7c087c3",
   876 => x"26487189",
   877 => x"5b5e0e4f",
   878 => x"4a710e5c",
   879 => x"724cd4ff",
   880 => x"87eac049",
   881 => x"029b4b70",
   882 => x"8bc187c2",
   883 => x"c848d0ff",
   884 => x"d5c178c5",
   885 => x"c649737c",
   886 => x"d1e3c131",
   887 => x"484abf97",
   888 => x"7c70b071",
   889 => x"c448d0ff",
   890 => x"fe487378",
   891 => x"5e0e87d5",
   892 => x"0e5d5c5b",
   893 => x"4c7186f8",
   894 => x"e4fb7ec0",
   895 => x"c04bc087",
   896 => x"bf97dbfa",
   897 => x"04a9c049",
   898 => x"f9fb87cf",
   899 => x"c083c187",
   900 => x"bf97dbfa",
   901 => x"f106ab49",
   902 => x"dbfac087",
   903 => x"cf02bf97",
   904 => x"87f2fa87",
   905 => x"02994970",
   906 => x"ecc087c6",
   907 => x"87f105a9",
   908 => x"e1fa4bc0",
   909 => x"fa4d7087",
   910 => x"a6c887dc",
   911 => x"87d6fa58",
   912 => x"83c14a70",
   913 => x"9749a4c8",
   914 => x"02ad4969",
   915 => x"ffc087c7",
   916 => x"e7c005ad",
   917 => x"49a4c987",
   918 => x"c4496997",
   919 => x"c702a966",
   920 => x"ffc04887",
   921 => x"87d405a8",
   922 => x"9749a4ca",
   923 => x"02aa4969",
   924 => x"ffc087c6",
   925 => x"87c405aa",
   926 => x"87d07ec1",
   927 => x"02adecc0",
   928 => x"fbc087c6",
   929 => x"87c405ad",
   930 => x"7ec14bc0",
   931 => x"e1fe026e",
   932 => x"87e9f987",
   933 => x"8ef84873",
   934 => x"0087e6fb",
   935 => x"5c5b5e0e",
   936 => x"711e0e5d",
   937 => x"4bd4ff4d",
   938 => x"e9c21e75",
   939 => x"fce649c8",
   940 => x"7086c487",
   941 => x"d8c30298",
   942 => x"d0e9c287",
   943 => x"49754cbf",
   944 => x"ff87f2fb",
   945 => x"c5c848d0",
   946 => x"7bd6c178",
   947 => x"a2754ac0",
   948 => x"c17b1149",
   949 => x"aab7cb82",
   950 => x"cc87f304",
   951 => x"7bffc34a",
   952 => x"e0c082c1",
   953 => x"f404aab7",
   954 => x"48d0ff87",
   955 => x"ffc378c4",
   956 => x"78c5c87b",
   957 => x"c17bd3c1",
   958 => x"7478c47b",
   959 => x"ffc1029c",
   960 => x"d2dcc287",
   961 => x"4dc0c87e",
   962 => x"acb7c08c",
   963 => x"c887c603",
   964 => x"c04da4c0",
   965 => x"adc0c84c",
   966 => x"c287dc05",
   967 => x"bf97c3e9",
   968 => x"0299d049",
   969 => x"1ec087d1",
   970 => x"49c8e9c2",
   971 => x"c487d3e8",
   972 => x"4a497086",
   973 => x"c287eec0",
   974 => x"c21ed2dc",
   975 => x"e849c8e9",
   976 => x"86c487c0",
   977 => x"ff4a4970",
   978 => x"c5c848d0",
   979 => x"7bd4c178",
   980 => x"7bbf976e",
   981 => x"80c1486e",
   982 => x"8dc17e70",
   983 => x"87f0ff05",
   984 => x"c448d0ff",
   985 => x"059a7278",
   986 => x"48c087c5",
   987 => x"c187e4c0",
   988 => x"c8e9c21e",
   989 => x"87f0e549",
   990 => x"9c7486c4",
   991 => x"87c1fe05",
   992 => x"c848d0ff",
   993 => x"d3c178c5",
   994 => x"c47bc07b",
   995 => x"c248c178",
   996 => x"2648c087",
   997 => x"4c264d26",
   998 => x"4f264b26",
   999 => x"5c5b5e0e",
  1000 => x"711e0e5d",
  1001 => x"4d4cc04b",
  1002 => x"e8c004ab",
  1003 => x"eef7c087",
  1004 => x"029d751e",
  1005 => x"4ac087c4",
  1006 => x"4ac187c2",
  1007 => x"dcec4972",
  1008 => x"7086c487",
  1009 => x"6e84c17e",
  1010 => x"7387c205",
  1011 => x"7385c14c",
  1012 => x"d8ff06ac",
  1013 => x"26486e87",
  1014 => x"0e87f9fe",
  1015 => x"0e5c5b5e",
  1016 => x"66cc4b71",
  1017 => x"4c87d802",
  1018 => x"028cf0c0",
  1019 => x"4a7487d8",
  1020 => x"d1028ac1",
  1021 => x"cd028a87",
  1022 => x"c9028a87",
  1023 => x"7387d987",
  1024 => x"87d8fa49",
  1025 => x"1e7487d2",
  1026 => x"d8c149c0",
  1027 => x"1e7487cb",
  1028 => x"d8c14973",
  1029 => x"86c887c3",
  1030 => x"0e87fbfd",
  1031 => x"5d5c5b5e",
  1032 => x"4c711e0e",
  1033 => x"c291de49",
  1034 => x"714df0e9",
  1035 => x"026d9785",
  1036 => x"c287dcc1",
  1037 => x"4abfdce9",
  1038 => x"49728274",
  1039 => x"7087ddfd",
  1040 => x"c0026e7e",
  1041 => x"e9c287f2",
  1042 => x"4a6e4be4",
  1043 => x"c1ff49cb",
  1044 => x"4b7487d6",
  1045 => x"e3c193cb",
  1046 => x"83c483e1",
  1047 => x"7bd3c2c1",
  1048 => x"c2c14974",
  1049 => x"7b7587cd",
  1050 => x"97d2e3c1",
  1051 => x"c21e49bf",
  1052 => x"fd49e4e9",
  1053 => x"86c487e5",
  1054 => x"c1c14974",
  1055 => x"49c087f5",
  1056 => x"87d4c3c1",
  1057 => x"48c4e9c2",
  1058 => x"49c178c0",
  1059 => x"2687c1dd",
  1060 => x"4c87c1fc",
  1061 => x"6964616f",
  1062 => x"2e2e676e",
  1063 => x"5e0e002e",
  1064 => x"710e5c5b",
  1065 => x"e9c24a4b",
  1066 => x"7282bfdc",
  1067 => x"87ecfb49",
  1068 => x"029c4c70",
  1069 => x"e74987c4",
  1070 => x"e9c287eb",
  1071 => x"78c048dc",
  1072 => x"cbdc49c1",
  1073 => x"87cefb87",
  1074 => x"5c5b5e0e",
  1075 => x"86f40e5d",
  1076 => x"4dd2dcc2",
  1077 => x"a6c44cc0",
  1078 => x"c278c048",
  1079 => x"49bfdce9",
  1080 => x"c106a9c0",
  1081 => x"dcc287c1",
  1082 => x"029848d2",
  1083 => x"c087f8c0",
  1084 => x"c81eeef7",
  1085 => x"87c70266",
  1086 => x"c048a6c4",
  1087 => x"c487c578",
  1088 => x"78c148a6",
  1089 => x"e74966c4",
  1090 => x"86c487d3",
  1091 => x"84c14d70",
  1092 => x"c14866c4",
  1093 => x"58a6c880",
  1094 => x"bfdce9c2",
  1095 => x"c603ac49",
  1096 => x"059d7587",
  1097 => x"c087c8ff",
  1098 => x"029d754c",
  1099 => x"c087e0c3",
  1100 => x"c81eeef7",
  1101 => x"87c70266",
  1102 => x"c048a6cc",
  1103 => x"cc87c578",
  1104 => x"78c148a6",
  1105 => x"e64966cc",
  1106 => x"86c487d3",
  1107 => x"026e7e70",
  1108 => x"6e87e9c2",
  1109 => x"9781cb49",
  1110 => x"99d04969",
  1111 => x"87d6c102",
  1112 => x"4adec2c1",
  1113 => x"91cb4974",
  1114 => x"81e1e3c1",
  1115 => x"81c87972",
  1116 => x"7451ffc3",
  1117 => x"c291de49",
  1118 => x"714df0e9",
  1119 => x"97c1c285",
  1120 => x"49a5c17d",
  1121 => x"c251e0c0",
  1122 => x"bf97e2e4",
  1123 => x"c187d202",
  1124 => x"4ba5c284",
  1125 => x"4ae2e4c2",
  1126 => x"fcfe49db",
  1127 => x"dbc187ca",
  1128 => x"49a5cd87",
  1129 => x"84c151c0",
  1130 => x"6e4ba5c2",
  1131 => x"fe49cb4a",
  1132 => x"c187f5fb",
  1133 => x"c0c187c6",
  1134 => x"49744adb",
  1135 => x"e3c191cb",
  1136 => x"797281e1",
  1137 => x"97e2e4c2",
  1138 => x"87d802bf",
  1139 => x"91de4974",
  1140 => x"e9c284c1",
  1141 => x"83714bf0",
  1142 => x"4ae2e4c2",
  1143 => x"fbfe49dd",
  1144 => x"87d887c6",
  1145 => x"93de4b74",
  1146 => x"83f0e9c2",
  1147 => x"c049a3cb",
  1148 => x"7384c151",
  1149 => x"49cb4a6e",
  1150 => x"87ecfafe",
  1151 => x"c14866c4",
  1152 => x"58a6c880",
  1153 => x"c003acc7",
  1154 => x"056e87c5",
  1155 => x"7487e0fc",
  1156 => x"f58ef448",
  1157 => x"731e87fe",
  1158 => x"494b711e",
  1159 => x"e3c191cb",
  1160 => x"a1c881e1",
  1161 => x"d1e3c14a",
  1162 => x"c9501248",
  1163 => x"fac04aa1",
  1164 => x"501248db",
  1165 => x"e3c181ca",
  1166 => x"501148d2",
  1167 => x"97d2e3c1",
  1168 => x"c01e49bf",
  1169 => x"87d3f649",
  1170 => x"48c4e9c2",
  1171 => x"49c178de",
  1172 => x"2687fdd5",
  1173 => x"1e87c1f5",
  1174 => x"cb494a71",
  1175 => x"e1e3c191",
  1176 => x"1181c881",
  1177 => x"c8e9c248",
  1178 => x"dce9c258",
  1179 => x"c178c048",
  1180 => x"87dcd549",
  1181 => x"c01e4f26",
  1182 => x"dbfbc049",
  1183 => x"1e4f2687",
  1184 => x"d2029971",
  1185 => x"f6e4c187",
  1186 => x"f750c048",
  1187 => x"d7c9c180",
  1188 => x"dae3c140",
  1189 => x"c187ce78",
  1190 => x"c148f2e4",
  1191 => x"fc78d3e3",
  1192 => x"f6c9c180",
  1193 => x"0e4f2678",
  1194 => x"0e5c5b5e",
  1195 => x"cb4a4c71",
  1196 => x"e1e3c192",
  1197 => x"49a2c882",
  1198 => x"974ba2c9",
  1199 => x"971e4b6b",
  1200 => x"ca1e4969",
  1201 => x"c0491282",
  1202 => x"c087d6e6",
  1203 => x"87c0d449",
  1204 => x"f8c04974",
  1205 => x"8ef887dd",
  1206 => x"1e87fbf2",
  1207 => x"4b711e73",
  1208 => x"87c3ff49",
  1209 => x"fefe4973",
  1210 => x"87ecf287",
  1211 => x"711e731e",
  1212 => x"4aa3c64b",
  1213 => x"c187db02",
  1214 => x"87d6028a",
  1215 => x"dac1028a",
  1216 => x"c0028a87",
  1217 => x"028a87fc",
  1218 => x"8a87e1c0",
  1219 => x"c187cb02",
  1220 => x"49c787db",
  1221 => x"c187c0fd",
  1222 => x"e9c287de",
  1223 => x"c102bfdc",
  1224 => x"c14887cb",
  1225 => x"e0e9c288",
  1226 => x"87c1c158",
  1227 => x"bfe0e9c2",
  1228 => x"87f9c002",
  1229 => x"bfdce9c2",
  1230 => x"c280c148",
  1231 => x"c058e0e9",
  1232 => x"e9c287eb",
  1233 => x"c649bfdc",
  1234 => x"e0e9c289",
  1235 => x"a9b7c059",
  1236 => x"c287da03",
  1237 => x"c048dce9",
  1238 => x"c287d278",
  1239 => x"02bfe0e9",
  1240 => x"e9c287cb",
  1241 => x"c648bfdc",
  1242 => x"e0e9c280",
  1243 => x"d149c058",
  1244 => x"497387de",
  1245 => x"87fbf5c0",
  1246 => x"0e87ddf0",
  1247 => x"0e5c5b5e",
  1248 => x"66cc4c71",
  1249 => x"cb4b741e",
  1250 => x"e1e3c193",
  1251 => x"4aa3c483",
  1252 => x"f4fe496a",
  1253 => x"c8c187e2",
  1254 => x"a3c87bd6",
  1255 => x"5166d449",
  1256 => x"d849a3c9",
  1257 => x"a3ca5166",
  1258 => x"5166dc49",
  1259 => x"87e6ef26",
  1260 => x"5c5b5e0e",
  1261 => x"d0ff0e5d",
  1262 => x"59a6d886",
  1263 => x"c048a6c4",
  1264 => x"c180c478",
  1265 => x"c47866c4",
  1266 => x"c478c180",
  1267 => x"c278c180",
  1268 => x"c148e0e9",
  1269 => x"c4e9c278",
  1270 => x"a8de48bf",
  1271 => x"f387cb05",
  1272 => x"497087e6",
  1273 => x"ce59a6c8",
  1274 => x"f4e387ee",
  1275 => x"87d6e487",
  1276 => x"7087e3e3",
  1277 => x"acfbc04c",
  1278 => x"87d0c102",
  1279 => x"c10566d4",
  1280 => x"1ec087c2",
  1281 => x"c11ec11e",
  1282 => x"c01ed4e5",
  1283 => x"87ebfd49",
  1284 => x"4a66d0c1",
  1285 => x"496a82c4",
  1286 => x"517481c7",
  1287 => x"1ed81ec1",
  1288 => x"81c8496a",
  1289 => x"d887f3e3",
  1290 => x"66c4c186",
  1291 => x"01a8c048",
  1292 => x"a6c487c7",
  1293 => x"ce78c148",
  1294 => x"66c4c187",
  1295 => x"cc88c148",
  1296 => x"87c358a6",
  1297 => x"cc87ffe2",
  1298 => x"78c248a6",
  1299 => x"cd029c74",
  1300 => x"66c487c2",
  1301 => x"66c8c148",
  1302 => x"f7cc03a8",
  1303 => x"48a6d887",
  1304 => x"80c478c0",
  1305 => x"ede178c0",
  1306 => x"c14c7087",
  1307 => x"c205acd0",
  1308 => x"66dc87d8",
  1309 => x"87d1e47e",
  1310 => x"e0c04970",
  1311 => x"d5e159a6",
  1312 => x"c04c7087",
  1313 => x"c105acec",
  1314 => x"66c487eb",
  1315 => x"c191cb49",
  1316 => x"c48166c0",
  1317 => x"4d6a4aa1",
  1318 => x"dc4aa1c8",
  1319 => x"c9c15266",
  1320 => x"f1e079d7",
  1321 => x"9c4c7087",
  1322 => x"c087d802",
  1323 => x"d202acfb",
  1324 => x"e0557487",
  1325 => x"4c7087e0",
  1326 => x"87c7029c",
  1327 => x"05acfbc0",
  1328 => x"c087eeff",
  1329 => x"c1c255e0",
  1330 => x"7d97c055",
  1331 => x"6e4966d4",
  1332 => x"87db05a9",
  1333 => x"c84866c4",
  1334 => x"ca04a866",
  1335 => x"4866c487",
  1336 => x"a6c880c1",
  1337 => x"c887c858",
  1338 => x"88c14866",
  1339 => x"ff58a6cc",
  1340 => x"7087e3df",
  1341 => x"acd0c14c",
  1342 => x"d087c805",
  1343 => x"80c14866",
  1344 => x"c158a6d4",
  1345 => x"fd02acd0",
  1346 => x"e0c087e8",
  1347 => x"66d448a6",
  1348 => x"4866dc78",
  1349 => x"a866e0c0",
  1350 => x"87cac905",
  1351 => x"48a6e4c0",
  1352 => x"747e78c0",
  1353 => x"88fbc048",
  1354 => x"58a6ecc0",
  1355 => x"c8029870",
  1356 => x"cb4887cf",
  1357 => x"a6ecc088",
  1358 => x"02987058",
  1359 => x"4887d2c1",
  1360 => x"ecc088c9",
  1361 => x"987058a6",
  1362 => x"87dbc302",
  1363 => x"c088c448",
  1364 => x"7058a6ec",
  1365 => x"87d00298",
  1366 => x"c088c148",
  1367 => x"7058a6ec",
  1368 => x"c2c30298",
  1369 => x"87d3c787",
  1370 => x"c048a6d8",
  1371 => x"ddff78f0",
  1372 => x"4c7087e4",
  1373 => x"02acecc0",
  1374 => x"dc87c3c0",
  1375 => x"ecc05ca6",
  1376 => x"87cd02ac",
  1377 => x"87ceddff",
  1378 => x"ecc04c70",
  1379 => x"f3ff05ac",
  1380 => x"acecc087",
  1381 => x"87c4c002",
  1382 => x"87fadcff",
  1383 => x"d41e66d8",
  1384 => x"d41e4966",
  1385 => x"c11e4966",
  1386 => x"d41ed4e5",
  1387 => x"caf74966",
  1388 => x"ca1ec087",
  1389 => x"4966dc1e",
  1390 => x"d8c191cb",
  1391 => x"a6d88166",
  1392 => x"78a1c448",
  1393 => x"49bf66d8",
  1394 => x"87ceddff",
  1395 => x"b7c086d8",
  1396 => x"c5c106a8",
  1397 => x"de1ec187",
  1398 => x"bf66c81e",
  1399 => x"f9dcff49",
  1400 => x"7086c887",
  1401 => x"08c04849",
  1402 => x"58a6dc88",
  1403 => x"06a8b7c0",
  1404 => x"d887e7c0",
  1405 => x"b7dd4866",
  1406 => x"87de03a8",
  1407 => x"d849bf6e",
  1408 => x"e0c08166",
  1409 => x"4966d851",
  1410 => x"bf6e81c1",
  1411 => x"51c1c281",
  1412 => x"c24966d8",
  1413 => x"81bf6e81",
  1414 => x"66cc51c0",
  1415 => x"d080c148",
  1416 => x"7ec158a6",
  1417 => x"ff87dac4",
  1418 => x"dc87dedd",
  1419 => x"ddff58a6",
  1420 => x"ecc087d7",
  1421 => x"ecc058a6",
  1422 => x"cac005a8",
  1423 => x"a6e8c087",
  1424 => x"7866d848",
  1425 => x"ff87c4c0",
  1426 => x"c487cbda",
  1427 => x"91cb4966",
  1428 => x"4866c0c1",
  1429 => x"7e708071",
  1430 => x"82c84a6e",
  1431 => x"81ca496e",
  1432 => x"c05166d8",
  1433 => x"c14966e8",
  1434 => x"8966d881",
  1435 => x"307148c1",
  1436 => x"89c14970",
  1437 => x"c27a9771",
  1438 => x"49bfcced",
  1439 => x"972966d8",
  1440 => x"71484a6a",
  1441 => x"a6f0c098",
  1442 => x"c4496e58",
  1443 => x"c04d6981",
  1444 => x"dc4866e0",
  1445 => x"c002a866",
  1446 => x"a6d887c8",
  1447 => x"c078c048",
  1448 => x"a6d887c5",
  1449 => x"d878c148",
  1450 => x"e0c01e66",
  1451 => x"ff49751e",
  1452 => x"c887e7d9",
  1453 => x"c04c7086",
  1454 => x"c106acb7",
  1455 => x"857487d4",
  1456 => x"7449e0c0",
  1457 => x"c14b7589",
  1458 => x"714acddf",
  1459 => x"87d8e7fe",
  1460 => x"e4c085c2",
  1461 => x"80c14866",
  1462 => x"58a6e8c0",
  1463 => x"4966ecc0",
  1464 => x"a97081c1",
  1465 => x"87c8c002",
  1466 => x"c048a6d8",
  1467 => x"87c5c078",
  1468 => x"c148a6d8",
  1469 => x"1e66d878",
  1470 => x"c049a4c2",
  1471 => x"887148e0",
  1472 => x"751e4970",
  1473 => x"d1d8ff49",
  1474 => x"c086c887",
  1475 => x"ff01a8b7",
  1476 => x"e4c087c0",
  1477 => x"d1c00266",
  1478 => x"c9496e87",
  1479 => x"66e4c081",
  1480 => x"c1486e51",
  1481 => x"c078e7ca",
  1482 => x"496e87cc",
  1483 => x"51c281c9",
  1484 => x"cbc1486e",
  1485 => x"7ec178db",
  1486 => x"ff87c6c0",
  1487 => x"7087c7d7",
  1488 => x"c0026e4c",
  1489 => x"66c487f5",
  1490 => x"a866c848",
  1491 => x"87cbc004",
  1492 => x"c14866c4",
  1493 => x"58a6c880",
  1494 => x"c887e0c0",
  1495 => x"88c14866",
  1496 => x"c058a6cc",
  1497 => x"c6c187d5",
  1498 => x"c8c005ac",
  1499 => x"4866cc87",
  1500 => x"a6d080c1",
  1501 => x"cdd6ff58",
  1502 => x"d04c7087",
  1503 => x"80c14866",
  1504 => x"7458a6d4",
  1505 => x"cbc0029c",
  1506 => x"4866c487",
  1507 => x"a866c8c1",
  1508 => x"87c9f304",
  1509 => x"87e5d5ff",
  1510 => x"c74866c4",
  1511 => x"e5c003a8",
  1512 => x"e0e9c287",
  1513 => x"c478c048",
  1514 => x"91cb4966",
  1515 => x"8166c0c1",
  1516 => x"6a4aa1c4",
  1517 => x"7952c04a",
  1518 => x"c14866c4",
  1519 => x"58a6c880",
  1520 => x"ff04a8c7",
  1521 => x"d0ff87db",
  1522 => x"c7dfff8e",
  1523 => x"00203a87",
  1524 => x"711e731e",
  1525 => x"c6029b4b",
  1526 => x"dce9c287",
  1527 => x"c778c048",
  1528 => x"dce9c21e",
  1529 => x"c11e49bf",
  1530 => x"c21ee1e3",
  1531 => x"49bfc4e9",
  1532 => x"cc87fdee",
  1533 => x"c4e9c286",
  1534 => x"c2ea49bf",
  1535 => x"029b7387",
  1536 => x"e3c187c8",
  1537 => x"e4c049e1",
  1538 => x"deff87fb",
  1539 => x"731e87ca",
  1540 => x"c14bc01e",
  1541 => x"c048d1e3",
  1542 => x"c4e5c150",
  1543 => x"d9ff49bf",
  1544 => x"987087fa",
  1545 => x"c187c405",
  1546 => x"734bf1e0",
  1547 => x"e7ddff48",
  1548 => x"4d4f5287",
  1549 => x"616f6c20",
  1550 => x"676e6964",
  1551 => x"69616620",
  1552 => x"0064656c",
  1553 => x"87ebc71e",
  1554 => x"c3fe49c1",
  1555 => x"cceafe87",
  1556 => x"02987087",
  1557 => x"f3fe87cd",
  1558 => x"987087c7",
  1559 => x"c187c402",
  1560 => x"c087c24a",
  1561 => x"059a724a",
  1562 => x"1ec087ce",
  1563 => x"49d8e2c1",
  1564 => x"87dfefc0",
  1565 => x"87fe86c4",
  1566 => x"87c7f9c0",
  1567 => x"e2c11ec0",
  1568 => x"efc049e3",
  1569 => x"1ec087cd",
  1570 => x"7087c3fe",
  1571 => x"c2efc049",
  1572 => x"87dec387",
  1573 => x"4f268ef8",
  1574 => x"66204453",
  1575 => x"656c6961",
  1576 => x"42002e64",
  1577 => x"69746f6f",
  1578 => x"2e2e676e",
  1579 => x"c01e002e",
  1580 => x"c087eee6",
  1581 => x"f687d2f2",
  1582 => x"1e4f2687",
  1583 => x"48dce9c2",
  1584 => x"e9c278c0",
  1585 => x"78c048c4",
  1586 => x"e187f9fd",
  1587 => x"2648c087",
  1588 => x"8000004f",
  1589 => x"69784520",
  1590 => x"20800074",
  1591 => x"6b636142",
  1592 => x"00125700",
  1593 => x"002a7000",
  1594 => x"00000000",
  1595 => x"00001257",
  1596 => x"00002a8e",
  1597 => x"57000000",
  1598 => x"ac000012",
  1599 => x"0000002a",
  1600 => x"12570000",
  1601 => x"2aca0000",
  1602 => x"00000000",
  1603 => x"00125700",
  1604 => x"002ae800",
  1605 => x"00000000",
  1606 => x"00001257",
  1607 => x"00002b06",
  1608 => x"57000000",
  1609 => x"24000012",
  1610 => x"0000002b",
  1611 => x"12570000",
  1612 => x"00000000",
  1613 => x"00000000",
  1614 => x"0012ec00",
  1615 => x"00000000",
  1616 => x"00000000",
  1617 => x"00001948",
  1618 => x"4553414c",
  1619 => x"30303552",
  1620 => x"004d4f52",
  1621 => x"64616f4c",
  1622 => x"002e2a20",
  1623 => x"48f0fe1e",
  1624 => x"09cd78c0",
  1625 => x"4f260979",
  1626 => x"f0fe1e1e",
  1627 => x"26487ebf",
  1628 => x"fe1e4f26",
  1629 => x"78c148f0",
  1630 => x"fe1e4f26",
  1631 => x"78c048f0",
  1632 => x"711e4f26",
  1633 => x"5252c04a",
  1634 => x"5e0e4f26",
  1635 => x"0e5d5c5b",
  1636 => x"4d7186f4",
  1637 => x"c17e6d97",
  1638 => x"6c974ca5",
  1639 => x"58a6c848",
  1640 => x"66c4486e",
  1641 => x"87c505a8",
  1642 => x"e6c048ff",
  1643 => x"87caff87",
  1644 => x"9749a5c2",
  1645 => x"a3714b6c",
  1646 => x"4b6b974b",
  1647 => x"6e7e6c97",
  1648 => x"c880c148",
  1649 => x"98c758a6",
  1650 => x"7058a6cc",
  1651 => x"e1fe7c97",
  1652 => x"f4487387",
  1653 => x"264d268e",
  1654 => x"264b264c",
  1655 => x"5b5e0e4f",
  1656 => x"86f40e5c",
  1657 => x"66d84c71",
  1658 => x"9affc34a",
  1659 => x"974ba4c2",
  1660 => x"a173496c",
  1661 => x"97517249",
  1662 => x"486e7e6c",
  1663 => x"a6c880c1",
  1664 => x"cc98c758",
  1665 => x"547058a6",
  1666 => x"caff8ef4",
  1667 => x"fd1e1e87",
  1668 => x"bfe087e8",
  1669 => x"e0c0494a",
  1670 => x"cb0299c0",
  1671 => x"c21e7287",
  1672 => x"fe49c2ed",
  1673 => x"86c487f7",
  1674 => x"7087fdfc",
  1675 => x"87c2fd7e",
  1676 => x"1e4f2626",
  1677 => x"49c2edc2",
  1678 => x"c187c7fd",
  1679 => x"fc49cde8",
  1680 => x"c8c487da",
  1681 => x"1e4f2687",
  1682 => x"c848d0ff",
  1683 => x"d4ff78e1",
  1684 => x"c478c548",
  1685 => x"87c30266",
  1686 => x"c878e0c3",
  1687 => x"87c60266",
  1688 => x"c348d4ff",
  1689 => x"d4ff78f0",
  1690 => x"ff787148",
  1691 => x"e1c848d0",
  1692 => x"78e0c078",
  1693 => x"5e0e4f26",
  1694 => x"710e5c5b",
  1695 => x"c2edc24c",
  1696 => x"87c6fc49",
  1697 => x"b7c04a70",
  1698 => x"e3c204aa",
  1699 => x"aae0c387",
  1700 => x"c187c905",
  1701 => x"c148c0ed",
  1702 => x"87d4c278",
  1703 => x"05aaf0c3",
  1704 => x"ecc187c9",
  1705 => x"78c148fc",
  1706 => x"c187f5c1",
  1707 => x"02bfc0ed",
  1708 => x"4b7287c7",
  1709 => x"c2b3c0c2",
  1710 => x"744b7287",
  1711 => x"87d1059c",
  1712 => x"bffcecc1",
  1713 => x"c0edc11e",
  1714 => x"49721ebf",
  1715 => x"c887f8fd",
  1716 => x"fcecc186",
  1717 => x"e0c002bf",
  1718 => x"c4497387",
  1719 => x"c19129b7",
  1720 => x"7381dcee",
  1721 => x"c29acf4a",
  1722 => x"7248c192",
  1723 => x"ff4a7030",
  1724 => x"694872ba",
  1725 => x"db797098",
  1726 => x"c4497387",
  1727 => x"c19129b7",
  1728 => x"7381dcee",
  1729 => x"c29acf4a",
  1730 => x"7248c392",
  1731 => x"484a7030",
  1732 => x"7970b069",
  1733 => x"48c0edc1",
  1734 => x"ecc178c0",
  1735 => x"78c048fc",
  1736 => x"49c2edc2",
  1737 => x"7087e3f9",
  1738 => x"aab7c04a",
  1739 => x"87ddfd03",
  1740 => x"87c248c0",
  1741 => x"4c264d26",
  1742 => x"4f264b26",
  1743 => x"00000000",
  1744 => x"00000000",
  1745 => x"494a711e",
  1746 => x"2687ebfc",
  1747 => x"4ac01e4f",
  1748 => x"91c44972",
  1749 => x"81dceec1",
  1750 => x"82c179c0",
  1751 => x"04aab7d0",
  1752 => x"4f2687ee",
  1753 => x"5c5b5e0e",
  1754 => x"4d710e5d",
  1755 => x"7587cbf8",
  1756 => x"2ab7c44a",
  1757 => x"dceec192",
  1758 => x"cf4c7582",
  1759 => x"6a94c29c",
  1760 => x"2b744b49",
  1761 => x"48c29bc3",
  1762 => x"4c703074",
  1763 => x"4874bcff",
  1764 => x"7a709871",
  1765 => x"7387dbf7",
  1766 => x"87d8fe48",
  1767 => x"00000000",
  1768 => x"00000000",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"48d0ff1e",
  1784 => x"7178e1c8",
  1785 => x"08d4ff48",
  1786 => x"1e4f2678",
  1787 => x"c848d0ff",
  1788 => x"487178e1",
  1789 => x"7808d4ff",
  1790 => x"ff4866c4",
  1791 => x"267808d4",
  1792 => x"4a711e4f",
  1793 => x"1e4966c4",
  1794 => x"deff4972",
  1795 => x"48d0ff87",
  1796 => x"2678e0c0",
  1797 => x"731e4f26",
  1798 => x"c84b711e",
  1799 => x"731e4966",
  1800 => x"a2e0c14a",
  1801 => x"87d9ff49",
  1802 => x"2687c426",
  1803 => x"264c264d",
  1804 => x"1e4f264b",
  1805 => x"c34ad4ff",
  1806 => x"d0ff7aff",
  1807 => x"78e1c848",
  1808 => x"edc27ade",
  1809 => x"497abfcc",
  1810 => x"7028c848",
  1811 => x"d048717a",
  1812 => x"717a7028",
  1813 => x"7028d848",
  1814 => x"48d0ff7a",
  1815 => x"2678e0c0",
  1816 => x"5b5e0e4f",
  1817 => x"710e5d5c",
  1818 => x"ccedc24c",
  1819 => x"744b4dbf",
  1820 => x"9b66d02b",
  1821 => x"66d483c1",
  1822 => x"87c204ab",
  1823 => x"4a744bc0",
  1824 => x"724966d0",
  1825 => x"75b9ff31",
  1826 => x"72487399",
  1827 => x"484a7030",
  1828 => x"edc2b071",
  1829 => x"dafe58d0",
  1830 => x"264d2687",
  1831 => x"264b264c",
  1832 => x"d0ff1e4f",
  1833 => x"78c9c848",
  1834 => x"d4ff4871",
  1835 => x"4f267808",
  1836 => x"494a711e",
  1837 => x"d0ff87eb",
  1838 => x"2678c848",
  1839 => x"1e731e4f",
  1840 => x"edc24b71",
  1841 => x"c302bfdc",
  1842 => x"87ebc287",
  1843 => x"c848d0ff",
  1844 => x"497378c9",
  1845 => x"ffb1e0c0",
  1846 => x"787148d4",
  1847 => x"48d0edc2",
  1848 => x"66c878c0",
  1849 => x"c387c502",
  1850 => x"87c249ff",
  1851 => x"edc249c0",
  1852 => x"66cc59d8",
  1853 => x"c587c602",
  1854 => x"c44ad5d5",
  1855 => x"ffffcf87",
  1856 => x"dcedc24a",
  1857 => x"dcedc25a",
  1858 => x"c478c148",
  1859 => x"264d2687",
  1860 => x"264b264c",
  1861 => x"5b5e0e4f",
  1862 => x"710e5d5c",
  1863 => x"d8edc24a",
  1864 => x"9a724cbf",
  1865 => x"4987cb02",
  1866 => x"f2c191c8",
  1867 => x"83714bf3",
  1868 => x"f6c187c4",
  1869 => x"4dc04bf3",
  1870 => x"99744913",
  1871 => x"bfd4edc2",
  1872 => x"48d4ffb9",
  1873 => x"b7c17871",
  1874 => x"b7c8852c",
  1875 => x"87e804ad",
  1876 => x"bfd0edc2",
  1877 => x"c280c848",
  1878 => x"fe58d4ed",
  1879 => x"731e87ef",
  1880 => x"134b711e",
  1881 => x"cb029a4a",
  1882 => x"fe497287",
  1883 => x"4a1387e7",
  1884 => x"87f5059a",
  1885 => x"1e87dafe",
  1886 => x"bfd0edc2",
  1887 => x"d0edc249",
  1888 => x"78a1c148",
  1889 => x"a9b7c0c4",
  1890 => x"ff87db03",
  1891 => x"edc248d4",
  1892 => x"c278bfd4",
  1893 => x"49bfd0ed",
  1894 => x"48d0edc2",
  1895 => x"c478a1c1",
  1896 => x"04a9b7c0",
  1897 => x"d0ff87e5",
  1898 => x"c278c848",
  1899 => x"c048dced",
  1900 => x"004f2678",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"5f5f0000",
  1904 => x"00000000",
  1905 => x"03000303",
  1906 => x"14000003",
  1907 => x"7f147f7f",
  1908 => x"0000147f",
  1909 => x"6b6b2e24",
  1910 => x"4c00123a",
  1911 => x"6c18366a",
  1912 => x"30003256",
  1913 => x"77594f7e",
  1914 => x"0040683a",
  1915 => x"03070400",
  1916 => x"00000000",
  1917 => x"633e1c00",
  1918 => x"00000041",
  1919 => x"3e634100",
  1920 => x"0800001c",
  1921 => x"1c1c3e2a",
  1922 => x"00082a3e",
  1923 => x"3e3e0808",
  1924 => x"00000808",
  1925 => x"60e08000",
  1926 => x"00000000",
  1927 => x"08080808",
  1928 => x"00000808",
  1929 => x"60600000",
  1930 => x"40000000",
  1931 => x"0c183060",
  1932 => x"00010306",
  1933 => x"4d597f3e",
  1934 => x"00003e7f",
  1935 => x"7f7f0604",
  1936 => x"00000000",
  1937 => x"59716342",
  1938 => x"0000464f",
  1939 => x"49496322",
  1940 => x"1800367f",
  1941 => x"7f13161c",
  1942 => x"0000107f",
  1943 => x"45456727",
  1944 => x"0000397d",
  1945 => x"494b7e3c",
  1946 => x"00003079",
  1947 => x"79710101",
  1948 => x"0000070f",
  1949 => x"49497f36",
  1950 => x"0000367f",
  1951 => x"69494f06",
  1952 => x"00001e3f",
  1953 => x"66660000",
  1954 => x"00000000",
  1955 => x"66e68000",
  1956 => x"00000000",
  1957 => x"14140808",
  1958 => x"00002222",
  1959 => x"14141414",
  1960 => x"00001414",
  1961 => x"14142222",
  1962 => x"00000808",
  1963 => x"59510302",
  1964 => x"3e00060f",
  1965 => x"555d417f",
  1966 => x"00001e1f",
  1967 => x"09097f7e",
  1968 => x"00007e7f",
  1969 => x"49497f7f",
  1970 => x"0000367f",
  1971 => x"41633e1c",
  1972 => x"00004141",
  1973 => x"63417f7f",
  1974 => x"00001c3e",
  1975 => x"49497f7f",
  1976 => x"00004141",
  1977 => x"09097f7f",
  1978 => x"00000101",
  1979 => x"49417f3e",
  1980 => x"00007a7b",
  1981 => x"08087f7f",
  1982 => x"00007f7f",
  1983 => x"7f7f4100",
  1984 => x"00000041",
  1985 => x"40406020",
  1986 => x"7f003f7f",
  1987 => x"361c087f",
  1988 => x"00004163",
  1989 => x"40407f7f",
  1990 => x"7f004040",
  1991 => x"060c067f",
  1992 => x"7f007f7f",
  1993 => x"180c067f",
  1994 => x"00007f7f",
  1995 => x"41417f3e",
  1996 => x"00003e7f",
  1997 => x"09097f7f",
  1998 => x"3e00060f",
  1999 => x"7f61417f",
  2000 => x"0000407e",
  2001 => x"19097f7f",
  2002 => x"0000667f",
  2003 => x"594d6f26",
  2004 => x"0000327b",
  2005 => x"7f7f0101",
  2006 => x"00000101",
  2007 => x"40407f3f",
  2008 => x"00003f7f",
  2009 => x"70703f0f",
  2010 => x"7f000f3f",
  2011 => x"3018307f",
  2012 => x"41007f7f",
  2013 => x"1c1c3663",
  2014 => x"01416336",
  2015 => x"7c7c0603",
  2016 => x"61010306",
  2017 => x"474d5971",
  2018 => x"00004143",
  2019 => x"417f7f00",
  2020 => x"01000041",
  2021 => x"180c0603",
  2022 => x"00406030",
  2023 => x"7f414100",
  2024 => x"0800007f",
  2025 => x"0603060c",
  2026 => x"8000080c",
  2027 => x"80808080",
  2028 => x"00008080",
  2029 => x"07030000",
  2030 => x"00000004",
  2031 => x"54547420",
  2032 => x"0000787c",
  2033 => x"44447f7f",
  2034 => x"0000387c",
  2035 => x"44447c38",
  2036 => x"00000044",
  2037 => x"44447c38",
  2038 => x"00007f7f",
  2039 => x"54547c38",
  2040 => x"0000185c",
  2041 => x"057f7e04",
  2042 => x"00000005",
  2043 => x"a4a4bc18",
  2044 => x"00007cfc",
  2045 => x"04047f7f",
  2046 => x"0000787c",
  2047 => x"7d3d0000",
  2048 => x"00000040",
  2049 => x"fd808080",
  2050 => x"0000007d",
  2051 => x"38107f7f",
  2052 => x"0000446c",
  2053 => x"7f3f0000",
  2054 => x"7c000040",
  2055 => x"0c180c7c",
  2056 => x"0000787c",
  2057 => x"04047c7c",
  2058 => x"0000787c",
  2059 => x"44447c38",
  2060 => x"0000387c",
  2061 => x"2424fcfc",
  2062 => x"0000183c",
  2063 => x"24243c18",
  2064 => x"0000fcfc",
  2065 => x"04047c7c",
  2066 => x"0000080c",
  2067 => x"54545c48",
  2068 => x"00002074",
  2069 => x"447f3f04",
  2070 => x"00000044",
  2071 => x"40407c3c",
  2072 => x"00007c7c",
  2073 => x"60603c1c",
  2074 => x"3c001c3c",
  2075 => x"6030607c",
  2076 => x"44003c7c",
  2077 => x"3810386c",
  2078 => x"0000446c",
  2079 => x"60e0bc1c",
  2080 => x"00001c3c",
  2081 => x"5c746444",
  2082 => x"0000444c",
  2083 => x"773e0808",
  2084 => x"00004141",
  2085 => x"7f7f0000",
  2086 => x"00000000",
  2087 => x"3e774141",
  2088 => x"02000808",
  2089 => x"02030101",
  2090 => x"7f000102",
  2091 => x"7f7f7f7f",
  2092 => x"08007f7f",
  2093 => x"3e1c1c08",
  2094 => x"7f7f7f3e",
  2095 => x"1c3e3e7f",
  2096 => x"0008081c",
  2097 => x"7c7c1810",
  2098 => x"00001018",
  2099 => x"7c7c3010",
  2100 => x"10001030",
  2101 => x"78606030",
  2102 => x"4200061e",
  2103 => x"3c183c66",
  2104 => x"78004266",
  2105 => x"c6c26a38",
  2106 => x"6000386c",
  2107 => x"00600000",
  2108 => x"0e006000",
  2109 => x"5d5c5b5e",
  2110 => x"4c711e0e",
  2111 => x"bfededc2",
  2112 => x"c04bc04d",
  2113 => x"02ab741e",
  2114 => x"a6c487c7",
  2115 => x"c578c048",
  2116 => x"48a6c487",
  2117 => x"66c478c1",
  2118 => x"ee49731e",
  2119 => x"86c887df",
  2120 => x"ef49e0c0",
  2121 => x"a5c487ef",
  2122 => x"f0496a4a",
  2123 => x"c6f187f0",
  2124 => x"c185cb87",
  2125 => x"abb7c883",
  2126 => x"87c7ff04",
  2127 => x"264d2626",
  2128 => x"264b264c",
  2129 => x"4a711e4f",
  2130 => x"5af1edc2",
  2131 => x"48f1edc2",
  2132 => x"fe4978c7",
  2133 => x"4f2687dd",
  2134 => x"711e731e",
  2135 => x"aab7c04a",
  2136 => x"c287d303",
  2137 => x"05bfe8d2",
  2138 => x"4bc187c4",
  2139 => x"4bc087c2",
  2140 => x"5becd2c2",
  2141 => x"d2c287c4",
  2142 => x"d2c25aec",
  2143 => x"c14abfe8",
  2144 => x"a2c0c19a",
  2145 => x"87e8ec49",
  2146 => x"d2c248fc",
  2147 => x"fe78bfe8",
  2148 => x"711e87ef",
  2149 => x"1e66c44a",
  2150 => x"f9e94972",
  2151 => x"4f262687",
  2152 => x"e8d2c21e",
  2153 => x"dbe649bf",
  2154 => x"e5edc287",
  2155 => x"78bfe848",
  2156 => x"48e1edc2",
  2157 => x"c278bfec",
  2158 => x"4abfe5ed",
  2159 => x"99ffc349",
  2160 => x"722ab7c8",
  2161 => x"c2b07148",
  2162 => x"2658eded",
  2163 => x"5b5e0e4f",
  2164 => x"710e5d5c",
  2165 => x"87c8ff4b",
  2166 => x"48e0edc2",
  2167 => x"497350c0",
  2168 => x"7087c1e6",
  2169 => x"9cc24c49",
  2170 => x"cb49eecb",
  2171 => x"497087c2",
  2172 => x"e0edc24d",
  2173 => x"c105bf97",
  2174 => x"66d087e2",
  2175 => x"e9edc249",
  2176 => x"d60599bf",
  2177 => x"4966d487",
  2178 => x"bfe1edc2",
  2179 => x"87cb0599",
  2180 => x"cfe54973",
  2181 => x"02987087",
  2182 => x"c187c1c1",
  2183 => x"87c0fe4c",
  2184 => x"d7ca4975",
  2185 => x"02987087",
  2186 => x"edc287c6",
  2187 => x"50c148e0",
  2188 => x"97e0edc2",
  2189 => x"e3c005bf",
  2190 => x"e9edc287",
  2191 => x"66d049bf",
  2192 => x"d6ff0599",
  2193 => x"e1edc287",
  2194 => x"66d449bf",
  2195 => x"caff0599",
  2196 => x"e4497387",
  2197 => x"987087ce",
  2198 => x"87fffe05",
  2199 => x"dcfb4874",
  2200 => x"5b5e0e87",
  2201 => x"f40e5d5c",
  2202 => x"4c4dc086",
  2203 => x"c47ebfec",
  2204 => x"edc248a6",
  2205 => x"c178bfed",
  2206 => x"c71ec01e",
  2207 => x"87cdfd49",
  2208 => x"987086c8",
  2209 => x"ff87cd02",
  2210 => x"87ccfb49",
  2211 => x"e349dac1",
  2212 => x"4dc187d2",
  2213 => x"97e0edc2",
  2214 => x"87c302bf",
  2215 => x"c287fbcf",
  2216 => x"4bbfe5ed",
  2217 => x"bfe8d2c2",
  2218 => x"87e9c005",
  2219 => x"e249fdc3",
  2220 => x"fac387f2",
  2221 => x"87ece249",
  2222 => x"ffc34973",
  2223 => x"c01e7199",
  2224 => x"87cefb49",
  2225 => x"b7c84973",
  2226 => x"c11e7129",
  2227 => x"87c2fb49",
  2228 => x"f9c586c8",
  2229 => x"e9edc287",
  2230 => x"029b4bbf",
  2231 => x"d2c287dd",
  2232 => x"c749bfe4",
  2233 => x"987087d6",
  2234 => x"c087c405",
  2235 => x"c287d24b",
  2236 => x"fbc649e0",
  2237 => x"e8d2c287",
  2238 => x"c287c658",
  2239 => x"c048e4d2",
  2240 => x"c2497378",
  2241 => x"87cd0599",
  2242 => x"e149ebc3",
  2243 => x"497087d6",
  2244 => x"c20299c2",
  2245 => x"734cfb87",
  2246 => x"0599c149",
  2247 => x"f4c387cd",
  2248 => x"87c0e149",
  2249 => x"99c24970",
  2250 => x"fa87c202",
  2251 => x"c849734c",
  2252 => x"87cd0599",
  2253 => x"e049f5c3",
  2254 => x"497087ea",
  2255 => x"d40299c2",
  2256 => x"f1edc287",
  2257 => x"87c902bf",
  2258 => x"c288c148",
  2259 => x"c258f5ed",
  2260 => x"c14cff87",
  2261 => x"c449734d",
  2262 => x"87cd0599",
  2263 => x"e049f2c3",
  2264 => x"497087c2",
  2265 => x"db0299c2",
  2266 => x"f1edc287",
  2267 => x"c7487ebf",
  2268 => x"cb03a8b7",
  2269 => x"c1486e87",
  2270 => x"f5edc280",
  2271 => x"87c2c058",
  2272 => x"4dc14cfe",
  2273 => x"ff49fdc3",
  2274 => x"7087d9df",
  2275 => x"0299c249",
  2276 => x"edc287d5",
  2277 => x"c002bff1",
  2278 => x"edc287c9",
  2279 => x"78c048f1",
  2280 => x"fd87c2c0",
  2281 => x"c34dc14c",
  2282 => x"deff49fa",
  2283 => x"497087f6",
  2284 => x"d90299c2",
  2285 => x"f1edc287",
  2286 => x"b7c748bf",
  2287 => x"c9c003a8",
  2288 => x"f1edc287",
  2289 => x"c078c748",
  2290 => x"4cfc87c2",
  2291 => x"b7c04dc1",
  2292 => x"d1c003ac",
  2293 => x"4a66c487",
  2294 => x"6a82d8c1",
  2295 => x"87c6c002",
  2296 => x"49744b6a",
  2297 => x"1ec00f73",
  2298 => x"c11ef0c3",
  2299 => x"dcf749da",
  2300 => x"7086c887",
  2301 => x"e2c00298",
  2302 => x"48a6c887",
  2303 => x"bff1edc2",
  2304 => x"4966c878",
  2305 => x"66c491cb",
  2306 => x"70807148",
  2307 => x"02bf6e7e",
  2308 => x"6e87c8c0",
  2309 => x"66c84bbf",
  2310 => x"750f7349",
  2311 => x"c8c0029d",
  2312 => x"f1edc287",
  2313 => x"caf349bf",
  2314 => x"ecd2c287",
  2315 => x"ddc002bf",
  2316 => x"c7c24987",
  2317 => x"02987087",
  2318 => x"c287d3c0",
  2319 => x"49bff1ed",
  2320 => x"c087f0f2",
  2321 => x"87d0f449",
  2322 => x"48ecd2c2",
  2323 => x"8ef478c0",
  2324 => x"0e87eaf3",
  2325 => x"5d5c5b5e",
  2326 => x"4c711e0e",
  2327 => x"bfededc2",
  2328 => x"a1cdc149",
  2329 => x"81d1c14d",
  2330 => x"9c747e69",
  2331 => x"c487cf02",
  2332 => x"7b744ba5",
  2333 => x"bfededc2",
  2334 => x"87c9f349",
  2335 => x"9c747b6e",
  2336 => x"c087c405",
  2337 => x"c187c24b",
  2338 => x"f349734b",
  2339 => x"66d487ca",
  2340 => x"4987c702",
  2341 => x"4a7087da",
  2342 => x"4ac087c2",
  2343 => x"5af0d2c2",
  2344 => x"87d9f226",
  2345 => x"00000000",
  2346 => x"00000000",
  2347 => x"00000000",
  2348 => x"ff4a711e",
  2349 => x"7249bfc8",
  2350 => x"4f2648a1",
  2351 => x"bfc8ff1e",
  2352 => x"c0c0fe89",
  2353 => x"a9c0c0c0",
  2354 => x"c087c401",
  2355 => x"c187c24a",
  2356 => x"2648724a",
  2357 => x"5b5e0e4f",
  2358 => x"710e5d5c",
  2359 => x"4cd4ff4b",
  2360 => x"c04866d0",
  2361 => x"ff49d678",
  2362 => x"c387f1db",
  2363 => x"496c7cff",
  2364 => x"7199ffc3",
  2365 => x"f0c3494d",
  2366 => x"a9e0c199",
  2367 => x"c387cb05",
  2368 => x"486c7cff",
  2369 => x"66d098c3",
  2370 => x"ffc37808",
  2371 => x"494a6c7c",
  2372 => x"ffc331c8",
  2373 => x"714a6c7c",
  2374 => x"c84972b2",
  2375 => x"7cffc331",
  2376 => x"b2714a6c",
  2377 => x"31c84972",
  2378 => x"6c7cffc3",
  2379 => x"ffb2714a",
  2380 => x"e0c048d0",
  2381 => x"029b7378",
  2382 => x"7b7287c2",
  2383 => x"4d264875",
  2384 => x"4b264c26",
  2385 => x"261e4f26",
  2386 => x"5b5e0e4f",
  2387 => x"86f80e5c",
  2388 => x"a6c81e76",
  2389 => x"87fdfd49",
  2390 => x"4b7086c4",
  2391 => x"a8c2486e",
  2392 => x"87f0c203",
  2393 => x"f0c34a73",
  2394 => x"aad0c19a",
  2395 => x"c187c702",
  2396 => x"c205aae0",
  2397 => x"497387de",
  2398 => x"c30299c8",
  2399 => x"87c6ff87",
  2400 => x"9cc34c73",
  2401 => x"c105acc2",
  2402 => x"66c487c2",
  2403 => x"7131c949",
  2404 => x"4a66c41e",
  2405 => x"edc292d4",
  2406 => x"817249f5",
  2407 => x"87c0d1fe",
  2408 => x"d8ff49d8",
  2409 => x"c0c887f6",
  2410 => x"d2dcc21e",
  2411 => x"fbecfd49",
  2412 => x"48d0ff87",
  2413 => x"c278e0c0",
  2414 => x"cc1ed2dc",
  2415 => x"92d44a66",
  2416 => x"49f5edc2",
  2417 => x"cffe8172",
  2418 => x"86cc87c7",
  2419 => x"c105acc1",
  2420 => x"66c487c2",
  2421 => x"7131c949",
  2422 => x"4a66c41e",
  2423 => x"edc292d4",
  2424 => x"817249f5",
  2425 => x"87f8cffe",
  2426 => x"1ed2dcc2",
  2427 => x"d44a66c8",
  2428 => x"f5edc292",
  2429 => x"fe817249",
  2430 => x"d787c7cd",
  2431 => x"dbd7ff49",
  2432 => x"1ec0c887",
  2433 => x"49d2dcc2",
  2434 => x"87f9eafd",
  2435 => x"d0ff86cc",
  2436 => x"78e0c048",
  2437 => x"e7fc8ef8",
  2438 => x"5b5e0e87",
  2439 => x"1e0e5d5c",
  2440 => x"d4ff4d71",
  2441 => x"7e66d44c",
  2442 => x"a8b7c348",
  2443 => x"c087c506",
  2444 => x"87e2c148",
  2445 => x"ddfe4975",
  2446 => x"1e7587fb",
  2447 => x"d44b66c4",
  2448 => x"f5edc293",
  2449 => x"fe497383",
  2450 => x"c887e2c8",
  2451 => x"ff4b6b83",
  2452 => x"e1c848d0",
  2453 => x"737cdd78",
  2454 => x"99ffc349",
  2455 => x"49737c71",
  2456 => x"c329b7c8",
  2457 => x"7c7199ff",
  2458 => x"b7d04973",
  2459 => x"99ffc329",
  2460 => x"49737c71",
  2461 => x"7129b7d8",
  2462 => x"7c7cc07c",
  2463 => x"7c7c7c7c",
  2464 => x"7c7c7c7c",
  2465 => x"e0c07c7c",
  2466 => x"1e66c478",
  2467 => x"d5ff49dc",
  2468 => x"86c887ef",
  2469 => x"fa264873",
  2470 => x"c21e87e4",
  2471 => x"49bfe8db",
  2472 => x"dbc2b9c1",
  2473 => x"d4ff59ec",
  2474 => x"78ffc348",
  2475 => x"c848d0ff",
  2476 => x"d4ff78e1",
  2477 => x"c478c148",
  2478 => x"ff787131",
  2479 => x"e0c048d0",
  2480 => x"1e4f2678",
  2481 => x"1edcdbc2",
  2482 => x"49c8e9c2",
  2483 => x"87ddc6fe",
  2484 => x"987086c4",
  2485 => x"ff87c302",
  2486 => x"4f2687c0",
  2487 => x"484b3531",
  2488 => x"2020205a",
  2489 => x"00474643",
  2490 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
