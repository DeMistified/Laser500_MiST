library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"00000040",
     1 => x"fd808080",
     2 => x"0000007d",
     3 => x"38107f7f",
     4 => x"0000446c",
     5 => x"7f3f0000",
     6 => x"7c000040",
     7 => x"0c180c7c",
     8 => x"0000787c",
     9 => x"04047c7c",
    10 => x"0000787c",
    11 => x"44447c38",
    12 => x"0000387c",
    13 => x"2424fcfc",
    14 => x"0000183c",
    15 => x"24243c18",
    16 => x"0000fcfc",
    17 => x"04047c7c",
    18 => x"0000080c",
    19 => x"54545c48",
    20 => x"00002074",
    21 => x"447f3f04",
    22 => x"00000044",
    23 => x"40407c3c",
    24 => x"00007c7c",
    25 => x"60603c1c",
    26 => x"3c001c3c",
    27 => x"6030607c",
    28 => x"44003c7c",
    29 => x"3810386c",
    30 => x"0000446c",
    31 => x"60e0bc1c",
    32 => x"00001c3c",
    33 => x"5c746444",
    34 => x"0000444c",
    35 => x"773e0808",
    36 => x"00004141",
    37 => x"7f7f0000",
    38 => x"00000000",
    39 => x"3e774141",
    40 => x"02000808",
    41 => x"02030101",
    42 => x"7f000102",
    43 => x"7f7f7f7f",
    44 => x"08007f7f",
    45 => x"3e1c1c08",
    46 => x"7f7f7f3e",
    47 => x"1c3e3e7f",
    48 => x"0008081c",
    49 => x"7c7c1810",
    50 => x"00001018",
    51 => x"7c7c3010",
    52 => x"10001030",
    53 => x"78606030",
    54 => x"4200061e",
    55 => x"3c183c66",
    56 => x"78004266",
    57 => x"c6c26a38",
    58 => x"6000386c",
    59 => x"00600000",
    60 => x"0e006000",
    61 => x"5d5c5b5e",
    62 => x"4c711e0e",
    63 => x"bfededc2",
    64 => x"c04bc04d",
    65 => x"02ab741e",
    66 => x"a6c487c7",
    67 => x"c578c048",
    68 => x"48a6c487",
    69 => x"66c478c1",
    70 => x"ee49731e",
    71 => x"86c887df",
    72 => x"ef49e0c0",
    73 => x"a5c487ef",
    74 => x"f0496a4a",
    75 => x"c6f187f0",
    76 => x"c185cb87",
    77 => x"abb7c883",
    78 => x"87c7ff04",
    79 => x"264d2626",
    80 => x"264b264c",
    81 => x"4a711e4f",
    82 => x"5af1edc2",
    83 => x"48f1edc2",
    84 => x"fe4978c7",
    85 => x"4f2687dd",
    86 => x"711e731e",
    87 => x"aab7c04a",
    88 => x"c287d303",
    89 => x"05bfe8d2",
    90 => x"4bc187c4",
    91 => x"4bc087c2",
    92 => x"5becd2c2",
    93 => x"d2c287c4",
    94 => x"d2c25aec",
    95 => x"c14abfe8",
    96 => x"a2c0c19a",
    97 => x"87e8ec49",
    98 => x"d2c248fc",
    99 => x"fe78bfe8",
   100 => x"711e87ef",
   101 => x"1e66c44a",
   102 => x"f9e94972",
   103 => x"4f262687",
   104 => x"e8d2c21e",
   105 => x"dbe649bf",
   106 => x"e5edc287",
   107 => x"78bfe848",
   108 => x"48e1edc2",
   109 => x"c278bfec",
   110 => x"4abfe5ed",
   111 => x"99ffc349",
   112 => x"722ab7c8",
   113 => x"c2b07148",
   114 => x"2658eded",
   115 => x"5b5e0e4f",
   116 => x"710e5d5c",
   117 => x"87c8ff4b",
   118 => x"48e0edc2",
   119 => x"497350c0",
   120 => x"7087c1e6",
   121 => x"9cc24c49",
   122 => x"cb49eecb",
   123 => x"497087c2",
   124 => x"e0edc24d",
   125 => x"c105bf97",
   126 => x"66d087e2",
   127 => x"e9edc249",
   128 => x"d60599bf",
   129 => x"4966d487",
   130 => x"bfe1edc2",
   131 => x"87cb0599",
   132 => x"cfe54973",
   133 => x"02987087",
   134 => x"c187c1c1",
   135 => x"87c0fe4c",
   136 => x"d7ca4975",
   137 => x"02987087",
   138 => x"edc287c6",
   139 => x"50c148e0",
   140 => x"97e0edc2",
   141 => x"e3c005bf",
   142 => x"e9edc287",
   143 => x"66d049bf",
   144 => x"d6ff0599",
   145 => x"e1edc287",
   146 => x"66d449bf",
   147 => x"caff0599",
   148 => x"e4497387",
   149 => x"987087ce",
   150 => x"87fffe05",
   151 => x"dcfb4874",
   152 => x"5b5e0e87",
   153 => x"f40e5d5c",
   154 => x"4c4dc086",
   155 => x"c47ebfec",
   156 => x"edc248a6",
   157 => x"c178bfed",
   158 => x"c71ec01e",
   159 => x"87cdfd49",
   160 => x"987086c8",
   161 => x"ff87cd02",
   162 => x"87ccfb49",
   163 => x"e349dac1",
   164 => x"4dc187d2",
   165 => x"97e0edc2",
   166 => x"87c302bf",
   167 => x"c287fbcf",
   168 => x"4bbfe5ed",
   169 => x"bfe8d2c2",
   170 => x"87e9c005",
   171 => x"e249fdc3",
   172 => x"fac387f2",
   173 => x"87ece249",
   174 => x"ffc34973",
   175 => x"c01e7199",
   176 => x"87cefb49",
   177 => x"b7c84973",
   178 => x"c11e7129",
   179 => x"87c2fb49",
   180 => x"f9c586c8",
   181 => x"e9edc287",
   182 => x"029b4bbf",
   183 => x"d2c287dd",
   184 => x"c749bfe4",
   185 => x"987087d6",
   186 => x"c087c405",
   187 => x"c287d24b",
   188 => x"fbc649e0",
   189 => x"e8d2c287",
   190 => x"c287c658",
   191 => x"c048e4d2",
   192 => x"c2497378",
   193 => x"87cd0599",
   194 => x"e149ebc3",
   195 => x"497087d6",
   196 => x"c20299c2",
   197 => x"734cfb87",
   198 => x"0599c149",
   199 => x"f4c387cd",
   200 => x"87c0e149",
   201 => x"99c24970",
   202 => x"fa87c202",
   203 => x"c849734c",
   204 => x"87cd0599",
   205 => x"e049f5c3",
   206 => x"497087ea",
   207 => x"d40299c2",
   208 => x"f1edc287",
   209 => x"87c902bf",
   210 => x"c288c148",
   211 => x"c258f5ed",
   212 => x"c14cff87",
   213 => x"c449734d",
   214 => x"87cd0599",
   215 => x"e049f2c3",
   216 => x"497087c2",
   217 => x"db0299c2",
   218 => x"f1edc287",
   219 => x"c7487ebf",
   220 => x"cb03a8b7",
   221 => x"c1486e87",
   222 => x"f5edc280",
   223 => x"87c2c058",
   224 => x"4dc14cfe",
   225 => x"ff49fdc3",
   226 => x"7087d9df",
   227 => x"0299c249",
   228 => x"edc287d5",
   229 => x"c002bff1",
   230 => x"edc287c9",
   231 => x"78c048f1",
   232 => x"fd87c2c0",
   233 => x"c34dc14c",
   234 => x"deff49fa",
   235 => x"497087f6",
   236 => x"d90299c2",
   237 => x"f1edc287",
   238 => x"b7c748bf",
   239 => x"c9c003a8",
   240 => x"f1edc287",
   241 => x"c078c748",
   242 => x"4cfc87c2",
   243 => x"b7c04dc1",
   244 => x"d1c003ac",
   245 => x"4a66c487",
   246 => x"6a82d8c1",
   247 => x"87c6c002",
   248 => x"49744b6a",
   249 => x"1ec00f73",
   250 => x"c11ef0c3",
   251 => x"dcf749da",
   252 => x"7086c887",
   253 => x"e2c00298",
   254 => x"48a6c887",
   255 => x"bff1edc2",
   256 => x"4966c878",
   257 => x"66c491cb",
   258 => x"70807148",
   259 => x"02bf6e7e",
   260 => x"6e87c8c0",
   261 => x"66c84bbf",
   262 => x"750f7349",
   263 => x"c8c0029d",
   264 => x"f1edc287",
   265 => x"caf349bf",
   266 => x"ecd2c287",
   267 => x"ddc002bf",
   268 => x"c7c24987",
   269 => x"02987087",
   270 => x"c287d3c0",
   271 => x"49bff1ed",
   272 => x"c087f0f2",
   273 => x"87d0f449",
   274 => x"48ecd2c2",
   275 => x"8ef478c0",
   276 => x"0e87eaf3",
   277 => x"5d5c5b5e",
   278 => x"4c711e0e",
   279 => x"bfededc2",
   280 => x"a1cdc149",
   281 => x"81d1c14d",
   282 => x"9c747e69",
   283 => x"c487cf02",
   284 => x"7b744ba5",
   285 => x"bfededc2",
   286 => x"87c9f349",
   287 => x"9c747b6e",
   288 => x"c087c405",
   289 => x"c187c24b",
   290 => x"f349734b",
   291 => x"66d487ca",
   292 => x"4987c702",
   293 => x"4a7087da",
   294 => x"4ac087c2",
   295 => x"5af0d2c2",
   296 => x"87d9f226",
   297 => x"00000000",
   298 => x"00000000",
   299 => x"00000000",
   300 => x"ff4a711e",
   301 => x"7249bfc8",
   302 => x"4f2648a1",
   303 => x"bfc8ff1e",
   304 => x"c0c0fe89",
   305 => x"a9c0c0c0",
   306 => x"c087c401",
   307 => x"c187c24a",
   308 => x"2648724a",
   309 => x"5b5e0e4f",
   310 => x"710e5d5c",
   311 => x"4cd4ff4b",
   312 => x"c04866d0",
   313 => x"ff49d678",
   314 => x"c387f1db",
   315 => x"496c7cff",
   316 => x"7199ffc3",
   317 => x"f0c3494d",
   318 => x"a9e0c199",
   319 => x"c387cb05",
   320 => x"486c7cff",
   321 => x"66d098c3",
   322 => x"ffc37808",
   323 => x"494a6c7c",
   324 => x"ffc331c8",
   325 => x"714a6c7c",
   326 => x"c84972b2",
   327 => x"7cffc331",
   328 => x"b2714a6c",
   329 => x"31c84972",
   330 => x"6c7cffc3",
   331 => x"ffb2714a",
   332 => x"e0c048d0",
   333 => x"029b7378",
   334 => x"7b7287c2",
   335 => x"4d264875",
   336 => x"4b264c26",
   337 => x"261e4f26",
   338 => x"5b5e0e4f",
   339 => x"86f80e5c",
   340 => x"a6c81e76",
   341 => x"87fdfd49",
   342 => x"4b7086c4",
   343 => x"a8c2486e",
   344 => x"87f0c203",
   345 => x"f0c34a73",
   346 => x"aad0c19a",
   347 => x"c187c702",
   348 => x"c205aae0",
   349 => x"497387de",
   350 => x"c30299c8",
   351 => x"87c6ff87",
   352 => x"9cc34c73",
   353 => x"c105acc2",
   354 => x"66c487c2",
   355 => x"7131c949",
   356 => x"4a66c41e",
   357 => x"edc292d4",
   358 => x"817249f5",
   359 => x"87c0d1fe",
   360 => x"d8ff49d8",
   361 => x"c0c887f6",
   362 => x"d2dcc21e",
   363 => x"fbecfd49",
   364 => x"48d0ff87",
   365 => x"c278e0c0",
   366 => x"cc1ed2dc",
   367 => x"92d44a66",
   368 => x"49f5edc2",
   369 => x"cffe8172",
   370 => x"86cc87c7",
   371 => x"c105acc1",
   372 => x"66c487c2",
   373 => x"7131c949",
   374 => x"4a66c41e",
   375 => x"edc292d4",
   376 => x"817249f5",
   377 => x"87f8cffe",
   378 => x"1ed2dcc2",
   379 => x"d44a66c8",
   380 => x"f5edc292",
   381 => x"fe817249",
   382 => x"d787c7cd",
   383 => x"dbd7ff49",
   384 => x"1ec0c887",
   385 => x"49d2dcc2",
   386 => x"87f9eafd",
   387 => x"d0ff86cc",
   388 => x"78e0c048",
   389 => x"e7fc8ef8",
   390 => x"5b5e0e87",
   391 => x"1e0e5d5c",
   392 => x"d4ff4d71",
   393 => x"7e66d44c",
   394 => x"a8b7c348",
   395 => x"c087c506",
   396 => x"87e2c148",
   397 => x"ddfe4975",
   398 => x"1e7587fb",
   399 => x"d44b66c4",
   400 => x"f5edc293",
   401 => x"fe497383",
   402 => x"c887e2c8",
   403 => x"ff4b6b83",
   404 => x"e1c848d0",
   405 => x"737cdd78",
   406 => x"99ffc349",
   407 => x"49737c71",
   408 => x"c329b7c8",
   409 => x"7c7199ff",
   410 => x"b7d04973",
   411 => x"99ffc329",
   412 => x"49737c71",
   413 => x"7129b7d8",
   414 => x"7c7cc07c",
   415 => x"7c7c7c7c",
   416 => x"7c7c7c7c",
   417 => x"e0c07c7c",
   418 => x"1e66c478",
   419 => x"d5ff49dc",
   420 => x"86c887ef",
   421 => x"fa264873",
   422 => x"c21e87e4",
   423 => x"49bfe8db",
   424 => x"dbc2b9c1",
   425 => x"d4ff59ec",
   426 => x"78ffc348",
   427 => x"c848d0ff",
   428 => x"d4ff78e1",
   429 => x"c478c148",
   430 => x"ff787131",
   431 => x"e0c048d0",
   432 => x"1e4f2678",
   433 => x"1edcdbc2",
   434 => x"49c8e9c2",
   435 => x"87ddc6fe",
   436 => x"987086c4",
   437 => x"ff87c302",
   438 => x"4f2687c0",
   439 => x"484b3531",
   440 => x"2020205a",
   441 => x"00474643",
   442 => x"00000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
