
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"e0",x"ee",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"e0",x"ee",x"c2"),
    14 => (x"48",x"ec",x"db",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"f0",x"e1"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"4a",x"71",x"1e",x"4f"),
    50 => (x"48",x"49",x"66",x"c4"),
    51 => (x"a6",x"c8",x"88",x"c1"),
    52 => (x"02",x"99",x"71",x"58"),
    53 => (x"48",x"12",x"87",x"d4"),
    54 => (x"78",x"08",x"d4",x"ff"),
    55 => (x"48",x"49",x"66",x"c4"),
    56 => (x"a6",x"c8",x"88",x"c1"),
    57 => (x"05",x"99",x"71",x"58"),
    58 => (x"4f",x"26",x"87",x"ec"),
    59 => (x"c4",x"4a",x"71",x"1e"),
    60 => (x"c1",x"48",x"49",x"66"),
    61 => (x"58",x"a6",x"c8",x"88"),
    62 => (x"d6",x"02",x"99",x"71"),
    63 => (x"48",x"d4",x"ff",x"87"),
    64 => (x"68",x"78",x"ff",x"c3"),
    65 => (x"49",x"66",x"c4",x"52"),
    66 => (x"c8",x"88",x"c1",x"48"),
    67 => (x"99",x"71",x"58",x"a6"),
    68 => (x"26",x"87",x"ea",x"05"),
    69 => (x"1e",x"73",x"1e",x"4f"),
    70 => (x"c3",x"4b",x"d4",x"ff"),
    71 => (x"4a",x"6b",x"7b",x"ff"),
    72 => (x"6b",x"7b",x"ff",x"c3"),
    73 => (x"72",x"32",x"c8",x"49"),
    74 => (x"7b",x"ff",x"c3",x"b1"),
    75 => (x"31",x"c8",x"4a",x"6b"),
    76 => (x"ff",x"c3",x"b2",x"71"),
    77 => (x"c8",x"49",x"6b",x"7b"),
    78 => (x"71",x"b1",x"72",x"32"),
    79 => (x"26",x"87",x"c4",x"48"),
    80 => (x"26",x"4c",x"26",x"4d"),
    81 => (x"0e",x"4f",x"26",x"4b"),
    82 => (x"5d",x"5c",x"5b",x"5e"),
    83 => (x"ff",x"4a",x"71",x"0e"),
    84 => (x"49",x"72",x"4c",x"d4"),
    85 => (x"71",x"99",x"ff",x"c3"),
    86 => (x"ec",x"db",x"c2",x"7c"),
    87 => (x"87",x"c8",x"05",x"bf"),
    88 => (x"c9",x"48",x"66",x"d0"),
    89 => (x"58",x"a6",x"d4",x"30"),
    90 => (x"d8",x"49",x"66",x"d0"),
    91 => (x"99",x"ff",x"c3",x"29"),
    92 => (x"66",x"d0",x"7c",x"71"),
    93 => (x"c3",x"29",x"d0",x"49"),
    94 => (x"7c",x"71",x"99",x"ff"),
    95 => (x"c8",x"49",x"66",x"d0"),
    96 => (x"99",x"ff",x"c3",x"29"),
    97 => (x"66",x"d0",x"7c",x"71"),
    98 => (x"99",x"ff",x"c3",x"49"),
    99 => (x"49",x"72",x"7c",x"71"),
   100 => (x"ff",x"c3",x"29",x"d0"),
   101 => (x"6c",x"7c",x"71",x"99"),
   102 => (x"ff",x"f0",x"c9",x"4b"),
   103 => (x"ab",x"ff",x"c3",x"4d"),
   104 => (x"c3",x"87",x"d0",x"05"),
   105 => (x"4b",x"6c",x"7c",x"ff"),
   106 => (x"c6",x"02",x"8d",x"c1"),
   107 => (x"ab",x"ff",x"c3",x"87"),
   108 => (x"73",x"87",x"f0",x"02"),
   109 => (x"87",x"c7",x"fe",x"48"),
   110 => (x"ff",x"49",x"c0",x"1e"),
   111 => (x"ff",x"c3",x"48",x"d4"),
   112 => (x"c3",x"81",x"c1",x"78"),
   113 => (x"04",x"a9",x"b7",x"c8"),
   114 => (x"4f",x"26",x"87",x"f1"),
   115 => (x"e7",x"1e",x"73",x"1e"),
   116 => (x"df",x"f8",x"c4",x"87"),
   117 => (x"c0",x"1e",x"c0",x"4b"),
   118 => (x"f7",x"c1",x"f0",x"ff"),
   119 => (x"87",x"e7",x"fd",x"49"),
   120 => (x"a8",x"c1",x"86",x"c4"),
   121 => (x"87",x"ea",x"c0",x"05"),
   122 => (x"c3",x"48",x"d4",x"ff"),
   123 => (x"c0",x"c1",x"78",x"ff"),
   124 => (x"c0",x"c0",x"c0",x"c0"),
   125 => (x"f0",x"e1",x"c0",x"1e"),
   126 => (x"fd",x"49",x"e9",x"c1"),
   127 => (x"86",x"c4",x"87",x"c9"),
   128 => (x"ca",x"05",x"98",x"70"),
   129 => (x"48",x"d4",x"ff",x"87"),
   130 => (x"c1",x"78",x"ff",x"c3"),
   131 => (x"fe",x"87",x"cb",x"48"),
   132 => (x"8b",x"c1",x"87",x"e6"),
   133 => (x"87",x"fd",x"fe",x"05"),
   134 => (x"e6",x"fc",x"48",x"c0"),
   135 => (x"1e",x"73",x"1e",x"87"),
   136 => (x"c3",x"48",x"d4",x"ff"),
   137 => (x"4b",x"d3",x"78",x"ff"),
   138 => (x"ff",x"c0",x"1e",x"c0"),
   139 => (x"49",x"c1",x"c1",x"f0"),
   140 => (x"c4",x"87",x"d4",x"fc"),
   141 => (x"05",x"98",x"70",x"86"),
   142 => (x"d4",x"ff",x"87",x"ca"),
   143 => (x"78",x"ff",x"c3",x"48"),
   144 => (x"87",x"cb",x"48",x"c1"),
   145 => (x"c1",x"87",x"f1",x"fd"),
   146 => (x"db",x"ff",x"05",x"8b"),
   147 => (x"fb",x"48",x"c0",x"87"),
   148 => (x"5e",x"0e",x"87",x"f1"),
   149 => (x"ff",x"0e",x"5c",x"5b"),
   150 => (x"db",x"fd",x"4c",x"d4"),
   151 => (x"1e",x"ea",x"c6",x"87"),
   152 => (x"c1",x"f0",x"e1",x"c0"),
   153 => (x"de",x"fb",x"49",x"c8"),
   154 => (x"c1",x"86",x"c4",x"87"),
   155 => (x"87",x"c8",x"02",x"a8"),
   156 => (x"c0",x"87",x"ea",x"fe"),
   157 => (x"87",x"e2",x"c1",x"48"),
   158 => (x"70",x"87",x"da",x"fa"),
   159 => (x"ff",x"ff",x"cf",x"49"),
   160 => (x"a9",x"ea",x"c6",x"99"),
   161 => (x"fe",x"87",x"c8",x"02"),
   162 => (x"48",x"c0",x"87",x"d3"),
   163 => (x"c3",x"87",x"cb",x"c1"),
   164 => (x"f1",x"c0",x"7c",x"ff"),
   165 => (x"87",x"f4",x"fc",x"4b"),
   166 => (x"c0",x"02",x"98",x"70"),
   167 => (x"1e",x"c0",x"87",x"eb"),
   168 => (x"c1",x"f0",x"ff",x"c0"),
   169 => (x"de",x"fa",x"49",x"fa"),
   170 => (x"70",x"86",x"c4",x"87"),
   171 => (x"87",x"d9",x"05",x"98"),
   172 => (x"6c",x"7c",x"ff",x"c3"),
   173 => (x"7c",x"ff",x"c3",x"49"),
   174 => (x"c1",x"7c",x"7c",x"7c"),
   175 => (x"c4",x"02",x"99",x"c0"),
   176 => (x"d5",x"48",x"c1",x"87"),
   177 => (x"d1",x"48",x"c0",x"87"),
   178 => (x"05",x"ab",x"c2",x"87"),
   179 => (x"48",x"c0",x"87",x"c4"),
   180 => (x"8b",x"c1",x"87",x"c8"),
   181 => (x"87",x"fd",x"fe",x"05"),
   182 => (x"e4",x"f9",x"48",x"c0"),
   183 => (x"1e",x"73",x"1e",x"87"),
   184 => (x"48",x"ec",x"db",x"c2"),
   185 => (x"4b",x"c7",x"78",x"c1"),
   186 => (x"c2",x"48",x"d0",x"ff"),
   187 => (x"87",x"c8",x"fb",x"78"),
   188 => (x"c3",x"48",x"d0",x"ff"),
   189 => (x"c0",x"1e",x"c0",x"78"),
   190 => (x"c0",x"c1",x"d0",x"e5"),
   191 => (x"87",x"c7",x"f9",x"49"),
   192 => (x"a8",x"c1",x"86",x"c4"),
   193 => (x"4b",x"87",x"c1",x"05"),
   194 => (x"c5",x"05",x"ab",x"c2"),
   195 => (x"c0",x"48",x"c0",x"87"),
   196 => (x"8b",x"c1",x"87",x"f9"),
   197 => (x"87",x"d0",x"ff",x"05"),
   198 => (x"c2",x"87",x"f7",x"fc"),
   199 => (x"70",x"58",x"f0",x"db"),
   200 => (x"87",x"cd",x"05",x"98"),
   201 => (x"ff",x"c0",x"1e",x"c1"),
   202 => (x"49",x"d0",x"c1",x"f0"),
   203 => (x"c4",x"87",x"d8",x"f8"),
   204 => (x"48",x"d4",x"ff",x"86"),
   205 => (x"c4",x"78",x"ff",x"c3"),
   206 => (x"db",x"c2",x"87",x"de"),
   207 => (x"d0",x"ff",x"58",x"f4"),
   208 => (x"ff",x"78",x"c2",x"48"),
   209 => (x"ff",x"c3",x"48",x"d4"),
   210 => (x"f7",x"48",x"c1",x"78"),
   211 => (x"5e",x"0e",x"87",x"f5"),
   212 => (x"0e",x"5d",x"5c",x"5b"),
   213 => (x"ff",x"c3",x"4a",x"71"),
   214 => (x"4c",x"d4",x"ff",x"4d"),
   215 => (x"d0",x"ff",x"7c",x"75"),
   216 => (x"78",x"c3",x"c4",x"48"),
   217 => (x"1e",x"72",x"7c",x"75"),
   218 => (x"c1",x"f0",x"ff",x"c0"),
   219 => (x"d6",x"f7",x"49",x"d8"),
   220 => (x"70",x"86",x"c4",x"87"),
   221 => (x"87",x"c5",x"02",x"98"),
   222 => (x"f0",x"c0",x"48",x"c1"),
   223 => (x"c3",x"7c",x"75",x"87"),
   224 => (x"c0",x"c8",x"7c",x"fe"),
   225 => (x"49",x"66",x"d4",x"1e"),
   226 => (x"c4",x"87",x"fa",x"f4"),
   227 => (x"75",x"7c",x"75",x"86"),
   228 => (x"d8",x"7c",x"75",x"7c"),
   229 => (x"75",x"4b",x"e0",x"da"),
   230 => (x"99",x"49",x"6c",x"7c"),
   231 => (x"c1",x"87",x"c5",x"05"),
   232 => (x"87",x"f3",x"05",x"8b"),
   233 => (x"d0",x"ff",x"7c",x"75"),
   234 => (x"c0",x"78",x"c2",x"48"),
   235 => (x"87",x"cf",x"f6",x"48"),
   236 => (x"5c",x"5b",x"5e",x"0e"),
   237 => (x"4b",x"71",x"0e",x"5d"),
   238 => (x"ee",x"c5",x"4c",x"c0"),
   239 => (x"ff",x"4a",x"df",x"cd"),
   240 => (x"ff",x"c3",x"48",x"d4"),
   241 => (x"c3",x"49",x"68",x"78"),
   242 => (x"c0",x"05",x"a9",x"fe"),
   243 => (x"4d",x"70",x"87",x"fd"),
   244 => (x"cc",x"02",x"9b",x"73"),
   245 => (x"1e",x"66",x"d0",x"87"),
   246 => (x"cf",x"f4",x"49",x"73"),
   247 => (x"d6",x"86",x"c4",x"87"),
   248 => (x"48",x"d0",x"ff",x"87"),
   249 => (x"c3",x"78",x"d1",x"c4"),
   250 => (x"66",x"d0",x"7d",x"ff"),
   251 => (x"d4",x"88",x"c1",x"48"),
   252 => (x"98",x"70",x"58",x"a6"),
   253 => (x"ff",x"87",x"f0",x"05"),
   254 => (x"ff",x"c3",x"48",x"d4"),
   255 => (x"9b",x"73",x"78",x"78"),
   256 => (x"ff",x"87",x"c5",x"05"),
   257 => (x"78",x"d0",x"48",x"d0"),
   258 => (x"c1",x"4c",x"4a",x"c1"),
   259 => (x"ee",x"fe",x"05",x"8a"),
   260 => (x"f4",x"48",x"74",x"87"),
   261 => (x"73",x"1e",x"87",x"e9"),
   262 => (x"c0",x"4a",x"71",x"1e"),
   263 => (x"48",x"d4",x"ff",x"4b"),
   264 => (x"ff",x"78",x"ff",x"c3"),
   265 => (x"c3",x"c4",x"48",x"d0"),
   266 => (x"48",x"d4",x"ff",x"78"),
   267 => (x"72",x"78",x"ff",x"c3"),
   268 => (x"f0",x"ff",x"c0",x"1e"),
   269 => (x"f4",x"49",x"d1",x"c1"),
   270 => (x"86",x"c4",x"87",x"cd"),
   271 => (x"d2",x"05",x"98",x"70"),
   272 => (x"1e",x"c0",x"c8",x"87"),
   273 => (x"fd",x"49",x"66",x"cc"),
   274 => (x"86",x"c4",x"87",x"e6"),
   275 => (x"d0",x"ff",x"4b",x"70"),
   276 => (x"73",x"78",x"c2",x"48"),
   277 => (x"87",x"eb",x"f3",x"48"),
   278 => (x"5c",x"5b",x"5e",x"0e"),
   279 => (x"1e",x"c0",x"0e",x"5d"),
   280 => (x"c1",x"f0",x"ff",x"c0"),
   281 => (x"de",x"f3",x"49",x"c9"),
   282 => (x"c2",x"1e",x"d2",x"87"),
   283 => (x"fc",x"49",x"f4",x"db"),
   284 => (x"86",x"c8",x"87",x"fe"),
   285 => (x"84",x"c1",x"4c",x"c0"),
   286 => (x"04",x"ac",x"b7",x"d2"),
   287 => (x"db",x"c2",x"87",x"f8"),
   288 => (x"49",x"bf",x"97",x"f4"),
   289 => (x"c1",x"99",x"c0",x"c3"),
   290 => (x"c0",x"05",x"a9",x"c0"),
   291 => (x"db",x"c2",x"87",x"e7"),
   292 => (x"49",x"bf",x"97",x"fb"),
   293 => (x"db",x"c2",x"31",x"d0"),
   294 => (x"4a",x"bf",x"97",x"fc"),
   295 => (x"b1",x"72",x"32",x"c8"),
   296 => (x"97",x"fd",x"db",x"c2"),
   297 => (x"71",x"b1",x"4a",x"bf"),
   298 => (x"ff",x"ff",x"cf",x"4c"),
   299 => (x"84",x"c1",x"9c",x"ff"),
   300 => (x"e7",x"c1",x"34",x"ca"),
   301 => (x"fd",x"db",x"c2",x"87"),
   302 => (x"c1",x"49",x"bf",x"97"),
   303 => (x"c2",x"99",x"c6",x"31"),
   304 => (x"bf",x"97",x"fe",x"db"),
   305 => (x"2a",x"b7",x"c7",x"4a"),
   306 => (x"db",x"c2",x"b1",x"72"),
   307 => (x"4a",x"bf",x"97",x"f9"),
   308 => (x"c2",x"9d",x"cf",x"4d"),
   309 => (x"bf",x"97",x"fa",x"db"),
   310 => (x"ca",x"9a",x"c3",x"4a"),
   311 => (x"fb",x"db",x"c2",x"32"),
   312 => (x"c2",x"4b",x"bf",x"97"),
   313 => (x"c2",x"b2",x"73",x"33"),
   314 => (x"bf",x"97",x"fc",x"db"),
   315 => (x"9b",x"c0",x"c3",x"4b"),
   316 => (x"73",x"2b",x"b7",x"c6"),
   317 => (x"c1",x"81",x"c2",x"b2"),
   318 => (x"70",x"30",x"71",x"48"),
   319 => (x"75",x"48",x"c1",x"49"),
   320 => (x"72",x"4d",x"70",x"30"),
   321 => (x"71",x"84",x"c1",x"4c"),
   322 => (x"b7",x"c0",x"c8",x"94"),
   323 => (x"87",x"cc",x"06",x"ad"),
   324 => (x"2d",x"b7",x"34",x"c1"),
   325 => (x"ad",x"b7",x"c0",x"c8"),
   326 => (x"87",x"f4",x"ff",x"01"),
   327 => (x"de",x"f0",x"48",x"74"),
   328 => (x"5b",x"5e",x"0e",x"87"),
   329 => (x"f8",x"0e",x"5d",x"5c"),
   330 => (x"da",x"e4",x"c2",x"86"),
   331 => (x"c2",x"78",x"c0",x"48"),
   332 => (x"c0",x"1e",x"d2",x"dc"),
   333 => (x"87",x"de",x"fb",x"49"),
   334 => (x"98",x"70",x"86",x"c4"),
   335 => (x"c0",x"87",x"c5",x"05"),
   336 => (x"87",x"ce",x"c9",x"48"),
   337 => (x"7e",x"c1",x"4d",x"c0"),
   338 => (x"bf",x"c0",x"f3",x"c0"),
   339 => (x"c8",x"dd",x"c2",x"49"),
   340 => (x"4b",x"c8",x"71",x"4a"),
   341 => (x"70",x"87",x"d3",x"ec"),
   342 => (x"87",x"c2",x"05",x"98"),
   343 => (x"f2",x"c0",x"7e",x"c0"),
   344 => (x"c2",x"49",x"bf",x"fc"),
   345 => (x"71",x"4a",x"e4",x"dd"),
   346 => (x"fd",x"eb",x"4b",x"c8"),
   347 => (x"05",x"98",x"70",x"87"),
   348 => (x"7e",x"c0",x"87",x"c2"),
   349 => (x"fd",x"c0",x"02",x"6e"),
   350 => (x"d8",x"e3",x"c2",x"87"),
   351 => (x"e4",x"c2",x"4d",x"bf"),
   352 => (x"7e",x"bf",x"9f",x"d0"),
   353 => (x"ea",x"d6",x"c5",x"48"),
   354 => (x"87",x"c7",x"05",x"a8"),
   355 => (x"bf",x"d8",x"e3",x"c2"),
   356 => (x"6e",x"87",x"ce",x"4d"),
   357 => (x"d5",x"e9",x"ca",x"48"),
   358 => (x"87",x"c5",x"02",x"a8"),
   359 => (x"f1",x"c7",x"48",x"c0"),
   360 => (x"d2",x"dc",x"c2",x"87"),
   361 => (x"f9",x"49",x"75",x"1e"),
   362 => (x"86",x"c4",x"87",x"ec"),
   363 => (x"c5",x"05",x"98",x"70"),
   364 => (x"c7",x"48",x"c0",x"87"),
   365 => (x"f2",x"c0",x"87",x"dc"),
   366 => (x"c2",x"49",x"bf",x"fc"),
   367 => (x"71",x"4a",x"e4",x"dd"),
   368 => (x"e5",x"ea",x"4b",x"c8"),
   369 => (x"05",x"98",x"70",x"87"),
   370 => (x"e4",x"c2",x"87",x"c8"),
   371 => (x"78",x"c1",x"48",x"da"),
   372 => (x"f3",x"c0",x"87",x"da"),
   373 => (x"c2",x"49",x"bf",x"c0"),
   374 => (x"71",x"4a",x"c8",x"dd"),
   375 => (x"c9",x"ea",x"4b",x"c8"),
   376 => (x"02",x"98",x"70",x"87"),
   377 => (x"c0",x"87",x"c5",x"c0"),
   378 => (x"87",x"e6",x"c6",x"48"),
   379 => (x"97",x"d0",x"e4",x"c2"),
   380 => (x"d5",x"c1",x"49",x"bf"),
   381 => (x"cd",x"c0",x"05",x"a9"),
   382 => (x"d1",x"e4",x"c2",x"87"),
   383 => (x"c2",x"49",x"bf",x"97"),
   384 => (x"c0",x"02",x"a9",x"ea"),
   385 => (x"48",x"c0",x"87",x"c5"),
   386 => (x"c2",x"87",x"c7",x"c6"),
   387 => (x"bf",x"97",x"d2",x"dc"),
   388 => (x"e9",x"c3",x"48",x"7e"),
   389 => (x"ce",x"c0",x"02",x"a8"),
   390 => (x"c3",x"48",x"6e",x"87"),
   391 => (x"c0",x"02",x"a8",x"eb"),
   392 => (x"48",x"c0",x"87",x"c5"),
   393 => (x"c2",x"87",x"eb",x"c5"),
   394 => (x"bf",x"97",x"dd",x"dc"),
   395 => (x"c0",x"05",x"99",x"49"),
   396 => (x"dc",x"c2",x"87",x"cc"),
   397 => (x"49",x"bf",x"97",x"de"),
   398 => (x"c0",x"02",x"a9",x"c2"),
   399 => (x"48",x"c0",x"87",x"c5"),
   400 => (x"c2",x"87",x"cf",x"c5"),
   401 => (x"bf",x"97",x"df",x"dc"),
   402 => (x"d6",x"e4",x"c2",x"48"),
   403 => (x"48",x"4c",x"70",x"58"),
   404 => (x"e4",x"c2",x"88",x"c1"),
   405 => (x"dc",x"c2",x"58",x"da"),
   406 => (x"49",x"bf",x"97",x"e0"),
   407 => (x"dc",x"c2",x"81",x"75"),
   408 => (x"4a",x"bf",x"97",x"e1"),
   409 => (x"a1",x"72",x"32",x"c8"),
   410 => (x"e7",x"e8",x"c2",x"7e"),
   411 => (x"c2",x"78",x"6e",x"48"),
   412 => (x"bf",x"97",x"e2",x"dc"),
   413 => (x"58",x"a6",x"c8",x"48"),
   414 => (x"bf",x"da",x"e4",x"c2"),
   415 => (x"87",x"d4",x"c2",x"02"),
   416 => (x"bf",x"fc",x"f2",x"c0"),
   417 => (x"e4",x"dd",x"c2",x"49"),
   418 => (x"4b",x"c8",x"71",x"4a"),
   419 => (x"70",x"87",x"db",x"e7"),
   420 => (x"c5",x"c0",x"02",x"98"),
   421 => (x"c3",x"48",x"c0",x"87"),
   422 => (x"e4",x"c2",x"87",x"f8"),
   423 => (x"c2",x"4c",x"bf",x"d2"),
   424 => (x"c2",x"5c",x"fb",x"e8"),
   425 => (x"bf",x"97",x"f7",x"dc"),
   426 => (x"c2",x"31",x"c8",x"49"),
   427 => (x"bf",x"97",x"f6",x"dc"),
   428 => (x"c2",x"49",x"a1",x"4a"),
   429 => (x"bf",x"97",x"f8",x"dc"),
   430 => (x"72",x"32",x"d0",x"4a"),
   431 => (x"dc",x"c2",x"49",x"a1"),
   432 => (x"4a",x"bf",x"97",x"f9"),
   433 => (x"a1",x"72",x"32",x"d8"),
   434 => (x"91",x"66",x"c4",x"49"),
   435 => (x"bf",x"e7",x"e8",x"c2"),
   436 => (x"ef",x"e8",x"c2",x"81"),
   437 => (x"ff",x"dc",x"c2",x"59"),
   438 => (x"c8",x"4a",x"bf",x"97"),
   439 => (x"fe",x"dc",x"c2",x"32"),
   440 => (x"a2",x"4b",x"bf",x"97"),
   441 => (x"c0",x"dd",x"c2",x"4a"),
   442 => (x"d0",x"4b",x"bf",x"97"),
   443 => (x"4a",x"a2",x"73",x"33"),
   444 => (x"97",x"c1",x"dd",x"c2"),
   445 => (x"9b",x"cf",x"4b",x"bf"),
   446 => (x"a2",x"73",x"33",x"d8"),
   447 => (x"f3",x"e8",x"c2",x"4a"),
   448 => (x"ef",x"e8",x"c2",x"5a"),
   449 => (x"8a",x"c2",x"4a",x"bf"),
   450 => (x"e8",x"c2",x"92",x"74"),
   451 => (x"a1",x"72",x"48",x"f3"),
   452 => (x"87",x"ca",x"c1",x"78"),
   453 => (x"97",x"e4",x"dc",x"c2"),
   454 => (x"31",x"c8",x"49",x"bf"),
   455 => (x"97",x"e3",x"dc",x"c2"),
   456 => (x"49",x"a1",x"4a",x"bf"),
   457 => (x"59",x"e2",x"e4",x"c2"),
   458 => (x"bf",x"de",x"e4",x"c2"),
   459 => (x"c7",x"31",x"c5",x"49"),
   460 => (x"29",x"c9",x"81",x"ff"),
   461 => (x"59",x"fb",x"e8",x"c2"),
   462 => (x"97",x"e9",x"dc",x"c2"),
   463 => (x"32",x"c8",x"4a",x"bf"),
   464 => (x"97",x"e8",x"dc",x"c2"),
   465 => (x"4a",x"a2",x"4b",x"bf"),
   466 => (x"6e",x"92",x"66",x"c4"),
   467 => (x"f7",x"e8",x"c2",x"82"),
   468 => (x"ef",x"e8",x"c2",x"5a"),
   469 => (x"c2",x"78",x"c0",x"48"),
   470 => (x"72",x"48",x"eb",x"e8"),
   471 => (x"e8",x"c2",x"78",x"a1"),
   472 => (x"e8",x"c2",x"48",x"fb"),
   473 => (x"c2",x"78",x"bf",x"ef"),
   474 => (x"c2",x"48",x"ff",x"e8"),
   475 => (x"78",x"bf",x"f3",x"e8"),
   476 => (x"bf",x"da",x"e4",x"c2"),
   477 => (x"87",x"c9",x"c0",x"02"),
   478 => (x"30",x"c4",x"48",x"74"),
   479 => (x"c9",x"c0",x"7e",x"70"),
   480 => (x"f7",x"e8",x"c2",x"87"),
   481 => (x"30",x"c4",x"48",x"bf"),
   482 => (x"e4",x"c2",x"7e",x"70"),
   483 => (x"78",x"6e",x"48",x"de"),
   484 => (x"8e",x"f8",x"48",x"c1"),
   485 => (x"4c",x"26",x"4d",x"26"),
   486 => (x"4f",x"26",x"4b",x"26"),
   487 => (x"5c",x"5b",x"5e",x"0e"),
   488 => (x"4a",x"71",x"0e",x"5d"),
   489 => (x"bf",x"da",x"e4",x"c2"),
   490 => (x"72",x"87",x"cb",x"02"),
   491 => (x"72",x"2b",x"c7",x"4b"),
   492 => (x"9c",x"ff",x"c1",x"4c"),
   493 => (x"4b",x"72",x"87",x"c9"),
   494 => (x"4c",x"72",x"2b",x"c8"),
   495 => (x"c2",x"9c",x"ff",x"c3"),
   496 => (x"83",x"bf",x"e7",x"e8"),
   497 => (x"bf",x"f8",x"f2",x"c0"),
   498 => (x"87",x"d9",x"02",x"ab"),
   499 => (x"5b",x"fc",x"f2",x"c0"),
   500 => (x"1e",x"d2",x"dc",x"c2"),
   501 => (x"fd",x"f0",x"49",x"73"),
   502 => (x"70",x"86",x"c4",x"87"),
   503 => (x"87",x"c5",x"05",x"98"),
   504 => (x"e6",x"c0",x"48",x"c0"),
   505 => (x"da",x"e4",x"c2",x"87"),
   506 => (x"87",x"d2",x"02",x"bf"),
   507 => (x"91",x"c4",x"49",x"74"),
   508 => (x"81",x"d2",x"dc",x"c2"),
   509 => (x"ff",x"cf",x"4d",x"69"),
   510 => (x"9d",x"ff",x"ff",x"ff"),
   511 => (x"49",x"74",x"87",x"cb"),
   512 => (x"dc",x"c2",x"91",x"c2"),
   513 => (x"69",x"9f",x"81",x"d2"),
   514 => (x"fe",x"48",x"75",x"4d"),
   515 => (x"5e",x"0e",x"87",x"c6"),
   516 => (x"0e",x"5d",x"5c",x"5b"),
   517 => (x"c0",x"4d",x"71",x"1e"),
   518 => (x"ca",x"49",x"c1",x"1e"),
   519 => (x"86",x"c4",x"87",x"ff"),
   520 => (x"02",x"9c",x"4c",x"70"),
   521 => (x"c2",x"87",x"c0",x"c1"),
   522 => (x"75",x"4a",x"e2",x"e4"),
   523 => (x"87",x"df",x"e0",x"49"),
   524 => (x"c0",x"02",x"98",x"70"),
   525 => (x"4a",x"74",x"87",x"f1"),
   526 => (x"4b",x"cb",x"49",x"75"),
   527 => (x"70",x"87",x"c5",x"e1"),
   528 => (x"e2",x"c0",x"02",x"98"),
   529 => (x"74",x"1e",x"c0",x"87"),
   530 => (x"87",x"c7",x"02",x"9c"),
   531 => (x"c0",x"48",x"a6",x"c4"),
   532 => (x"c4",x"87",x"c5",x"78"),
   533 => (x"78",x"c1",x"48",x"a6"),
   534 => (x"c9",x"49",x"66",x"c4"),
   535 => (x"86",x"c4",x"87",x"ff"),
   536 => (x"05",x"9c",x"4c",x"70"),
   537 => (x"74",x"87",x"c0",x"ff"),
   538 => (x"e7",x"fc",x"26",x"48"),
   539 => (x"5b",x"5e",x"0e",x"87"),
   540 => (x"1e",x"0e",x"5d",x"5c"),
   541 => (x"05",x"9b",x"4b",x"71"),
   542 => (x"48",x"c0",x"87",x"c5"),
   543 => (x"c8",x"87",x"e5",x"c1"),
   544 => (x"7d",x"c0",x"4d",x"a3"),
   545 => (x"c7",x"02",x"66",x"d4"),
   546 => (x"97",x"66",x"d4",x"87"),
   547 => (x"87",x"c5",x"05",x"bf"),
   548 => (x"cf",x"c1",x"48",x"c0"),
   549 => (x"49",x"66",x"d4",x"87"),
   550 => (x"70",x"87",x"f3",x"fd"),
   551 => (x"c1",x"02",x"9c",x"4c"),
   552 => (x"a4",x"dc",x"87",x"c0"),
   553 => (x"da",x"7d",x"69",x"49"),
   554 => (x"a3",x"c4",x"49",x"a4"),
   555 => (x"7a",x"69",x"9f",x"4a"),
   556 => (x"bf",x"da",x"e4",x"c2"),
   557 => (x"d4",x"87",x"d2",x"02"),
   558 => (x"69",x"9f",x"49",x"a4"),
   559 => (x"ff",x"ff",x"c0",x"49"),
   560 => (x"d0",x"48",x"71",x"99"),
   561 => (x"c2",x"7e",x"70",x"30"),
   562 => (x"6e",x"7e",x"c0",x"87"),
   563 => (x"80",x"6a",x"48",x"49"),
   564 => (x"7b",x"c0",x"7a",x"70"),
   565 => (x"6a",x"49",x"a3",x"cc"),
   566 => (x"49",x"a3",x"d0",x"79"),
   567 => (x"48",x"c1",x"79",x"c0"),
   568 => (x"48",x"c0",x"87",x"c2"),
   569 => (x"87",x"ec",x"fa",x"26"),
   570 => (x"5c",x"5b",x"5e",x"0e"),
   571 => (x"4c",x"71",x"0e",x"5d"),
   572 => (x"ca",x"c1",x"02",x"9c"),
   573 => (x"49",x"a4",x"c8",x"87"),
   574 => (x"c2",x"c1",x"02",x"69"),
   575 => (x"4a",x"66",x"d0",x"87"),
   576 => (x"d4",x"82",x"49",x"6c"),
   577 => (x"66",x"d0",x"5a",x"a6"),
   578 => (x"e4",x"c2",x"b9",x"4d"),
   579 => (x"ff",x"4a",x"bf",x"d6"),
   580 => (x"71",x"99",x"72",x"ba"),
   581 => (x"e4",x"c0",x"02",x"99"),
   582 => (x"4b",x"a4",x"c4",x"87"),
   583 => (x"fb",x"f9",x"49",x"6b"),
   584 => (x"c2",x"7b",x"70",x"87"),
   585 => (x"49",x"bf",x"d2",x"e4"),
   586 => (x"7c",x"71",x"81",x"6c"),
   587 => (x"e4",x"c2",x"b9",x"75"),
   588 => (x"ff",x"4a",x"bf",x"d6"),
   589 => (x"71",x"99",x"72",x"ba"),
   590 => (x"dc",x"ff",x"05",x"99"),
   591 => (x"f9",x"7c",x"75",x"87"),
   592 => (x"73",x"1e",x"87",x"d2"),
   593 => (x"9b",x"4b",x"71",x"1e"),
   594 => (x"c8",x"87",x"c7",x"02"),
   595 => (x"05",x"69",x"49",x"a3"),
   596 => (x"48",x"c0",x"87",x"c5"),
   597 => (x"c2",x"87",x"f7",x"c0"),
   598 => (x"4a",x"bf",x"eb",x"e8"),
   599 => (x"69",x"49",x"a3",x"c4"),
   600 => (x"c2",x"89",x"c2",x"49"),
   601 => (x"91",x"bf",x"d2",x"e4"),
   602 => (x"c2",x"4a",x"a2",x"71"),
   603 => (x"49",x"bf",x"d6",x"e4"),
   604 => (x"a2",x"71",x"99",x"6b"),
   605 => (x"fc",x"f2",x"c0",x"4a"),
   606 => (x"1e",x"66",x"c8",x"5a"),
   607 => (x"d5",x"ea",x"49",x"72"),
   608 => (x"70",x"86",x"c4",x"87"),
   609 => (x"87",x"c4",x"05",x"98"),
   610 => (x"87",x"c2",x"48",x"c0"),
   611 => (x"c7",x"f8",x"48",x"c1"),
   612 => (x"1e",x"73",x"1e",x"87"),
   613 => (x"02",x"9b",x"4b",x"71"),
   614 => (x"a3",x"c8",x"87",x"c7"),
   615 => (x"c5",x"05",x"69",x"49"),
   616 => (x"c0",x"48",x"c0",x"87"),
   617 => (x"e8",x"c2",x"87",x"f7"),
   618 => (x"c4",x"4a",x"bf",x"eb"),
   619 => (x"49",x"69",x"49",x"a3"),
   620 => (x"e4",x"c2",x"89",x"c2"),
   621 => (x"71",x"91",x"bf",x"d2"),
   622 => (x"e4",x"c2",x"4a",x"a2"),
   623 => (x"6b",x"49",x"bf",x"d6"),
   624 => (x"4a",x"a2",x"71",x"99"),
   625 => (x"5a",x"fc",x"f2",x"c0"),
   626 => (x"72",x"1e",x"66",x"c8"),
   627 => (x"87",x"fe",x"e5",x"49"),
   628 => (x"98",x"70",x"86",x"c4"),
   629 => (x"c0",x"87",x"c4",x"05"),
   630 => (x"c1",x"87",x"c2",x"48"),
   631 => (x"87",x"f8",x"f6",x"48"),
   632 => (x"5c",x"5b",x"5e",x"0e"),
   633 => (x"71",x"1e",x"0e",x"5d"),
   634 => (x"4c",x"66",x"d4",x"4b"),
   635 => (x"9b",x"73",x"2c",x"c9"),
   636 => (x"87",x"cf",x"c1",x"02"),
   637 => (x"69",x"49",x"a3",x"c8"),
   638 => (x"87",x"c7",x"c1",x"02"),
   639 => (x"d4",x"4d",x"a3",x"d0"),
   640 => (x"e4",x"c2",x"7d",x"66"),
   641 => (x"ff",x"49",x"bf",x"d6"),
   642 => (x"99",x"4a",x"6b",x"b9"),
   643 => (x"03",x"ac",x"71",x"7e"),
   644 => (x"7b",x"c0",x"87",x"cd"),
   645 => (x"4a",x"a3",x"cc",x"7d"),
   646 => (x"6a",x"49",x"a3",x"c4"),
   647 => (x"72",x"87",x"c2",x"79"),
   648 => (x"02",x"9c",x"74",x"8c"),
   649 => (x"1e",x"49",x"87",x"dd"),
   650 => (x"fb",x"fa",x"49",x"73"),
   651 => (x"d4",x"86",x"c4",x"87"),
   652 => (x"ff",x"c7",x"49",x"66"),
   653 => (x"87",x"cb",x"02",x"99"),
   654 => (x"1e",x"d2",x"dc",x"c2"),
   655 => (x"c1",x"fc",x"49",x"73"),
   656 => (x"26",x"86",x"c4",x"87"),
   657 => (x"1e",x"87",x"cd",x"f5"),
   658 => (x"4b",x"71",x"1e",x"73"),
   659 => (x"e4",x"c0",x"02",x"9b"),
   660 => (x"ff",x"e8",x"c2",x"87"),
   661 => (x"c2",x"4a",x"73",x"5b"),
   662 => (x"d2",x"e4",x"c2",x"8a"),
   663 => (x"c2",x"92",x"49",x"bf"),
   664 => (x"48",x"bf",x"eb",x"e8"),
   665 => (x"e9",x"c2",x"80",x"72"),
   666 => (x"48",x"71",x"58",x"c3"),
   667 => (x"e4",x"c2",x"30",x"c4"),
   668 => (x"ed",x"c0",x"58",x"e2"),
   669 => (x"fb",x"e8",x"c2",x"87"),
   670 => (x"ef",x"e8",x"c2",x"48"),
   671 => (x"e8",x"c2",x"78",x"bf"),
   672 => (x"e8",x"c2",x"48",x"ff"),
   673 => (x"c2",x"78",x"bf",x"f3"),
   674 => (x"02",x"bf",x"da",x"e4"),
   675 => (x"e4",x"c2",x"87",x"c9"),
   676 => (x"c4",x"49",x"bf",x"d2"),
   677 => (x"c2",x"87",x"c7",x"31"),
   678 => (x"49",x"bf",x"f7",x"e8"),
   679 => (x"e4",x"c2",x"31",x"c4"),
   680 => (x"f3",x"f3",x"59",x"e2"),
   681 => (x"5b",x"5e",x"0e",x"87"),
   682 => (x"4a",x"71",x"0e",x"5c"),
   683 => (x"9a",x"72",x"4b",x"c0"),
   684 => (x"87",x"e1",x"c0",x"02"),
   685 => (x"9f",x"49",x"a2",x"da"),
   686 => (x"e4",x"c2",x"4b",x"69"),
   687 => (x"cf",x"02",x"bf",x"da"),
   688 => (x"49",x"a2",x"d4",x"87"),
   689 => (x"4c",x"49",x"69",x"9f"),
   690 => (x"9c",x"ff",x"ff",x"c0"),
   691 => (x"87",x"c2",x"34",x"d0"),
   692 => (x"49",x"74",x"4c",x"c0"),
   693 => (x"fd",x"49",x"73",x"b3"),
   694 => (x"f9",x"f2",x"87",x"ed"),
   695 => (x"5b",x"5e",x"0e",x"87"),
   696 => (x"f4",x"0e",x"5d",x"5c"),
   697 => (x"c0",x"4a",x"71",x"86"),
   698 => (x"02",x"9a",x"72",x"7e"),
   699 => (x"dc",x"c2",x"87",x"d8"),
   700 => (x"78",x"c0",x"48",x"ce"),
   701 => (x"48",x"c6",x"dc",x"c2"),
   702 => (x"bf",x"ff",x"e8",x"c2"),
   703 => (x"ca",x"dc",x"c2",x"78"),
   704 => (x"fb",x"e8",x"c2",x"48"),
   705 => (x"e4",x"c2",x"78",x"bf"),
   706 => (x"50",x"c0",x"48",x"ef"),
   707 => (x"bf",x"de",x"e4",x"c2"),
   708 => (x"ce",x"dc",x"c2",x"49"),
   709 => (x"aa",x"71",x"4a",x"bf"),
   710 => (x"87",x"c9",x"c4",x"03"),
   711 => (x"99",x"cf",x"49",x"72"),
   712 => (x"87",x"e9",x"c0",x"05"),
   713 => (x"48",x"f8",x"f2",x"c0"),
   714 => (x"bf",x"c6",x"dc",x"c2"),
   715 => (x"d2",x"dc",x"c2",x"78"),
   716 => (x"c6",x"dc",x"c2",x"1e"),
   717 => (x"dc",x"c2",x"49",x"bf"),
   718 => (x"a1",x"c1",x"48",x"c6"),
   719 => (x"d5",x"e3",x"71",x"78"),
   720 => (x"c0",x"86",x"c4",x"87"),
   721 => (x"c2",x"48",x"f4",x"f2"),
   722 => (x"cc",x"78",x"d2",x"dc"),
   723 => (x"f4",x"f2",x"c0",x"87"),
   724 => (x"e0",x"c0",x"48",x"bf"),
   725 => (x"f8",x"f2",x"c0",x"80"),
   726 => (x"ce",x"dc",x"c2",x"58"),
   727 => (x"80",x"c1",x"48",x"bf"),
   728 => (x"58",x"d2",x"dc",x"c2"),
   729 => (x"00",x"0c",x"b4",x"27"),
   730 => (x"bf",x"97",x"bf",x"00"),
   731 => (x"c2",x"02",x"9d",x"4d"),
   732 => (x"e5",x"c3",x"87",x"e3"),
   733 => (x"dc",x"c2",x"02",x"ad"),
   734 => (x"f4",x"f2",x"c0",x"87"),
   735 => (x"a3",x"cb",x"4b",x"bf"),
   736 => (x"cf",x"4c",x"11",x"49"),
   737 => (x"d2",x"c1",x"05",x"ac"),
   738 => (x"df",x"49",x"75",x"87"),
   739 => (x"cd",x"89",x"c1",x"99"),
   740 => (x"e2",x"e4",x"c2",x"91"),
   741 => (x"4a",x"a3",x"c1",x"81"),
   742 => (x"a3",x"c3",x"51",x"12"),
   743 => (x"c5",x"51",x"12",x"4a"),
   744 => (x"51",x"12",x"4a",x"a3"),
   745 => (x"12",x"4a",x"a3",x"c7"),
   746 => (x"4a",x"a3",x"c9",x"51"),
   747 => (x"a3",x"ce",x"51",x"12"),
   748 => (x"d0",x"51",x"12",x"4a"),
   749 => (x"51",x"12",x"4a",x"a3"),
   750 => (x"12",x"4a",x"a3",x"d2"),
   751 => (x"4a",x"a3",x"d4",x"51"),
   752 => (x"a3",x"d6",x"51",x"12"),
   753 => (x"d8",x"51",x"12",x"4a"),
   754 => (x"51",x"12",x"4a",x"a3"),
   755 => (x"12",x"4a",x"a3",x"dc"),
   756 => (x"4a",x"a3",x"de",x"51"),
   757 => (x"7e",x"c1",x"51",x"12"),
   758 => (x"74",x"87",x"fa",x"c0"),
   759 => (x"05",x"99",x"c8",x"49"),
   760 => (x"74",x"87",x"eb",x"c0"),
   761 => (x"05",x"99",x"d0",x"49"),
   762 => (x"66",x"dc",x"87",x"d1"),
   763 => (x"87",x"cb",x"c0",x"02"),
   764 => (x"66",x"dc",x"49",x"73"),
   765 => (x"02",x"98",x"70",x"0f"),
   766 => (x"6e",x"87",x"d3",x"c0"),
   767 => (x"87",x"c6",x"c0",x"05"),
   768 => (x"48",x"e2",x"e4",x"c2"),
   769 => (x"f2",x"c0",x"50",x"c0"),
   770 => (x"c2",x"48",x"bf",x"f4"),
   771 => (x"e4",x"c2",x"87",x"e1"),
   772 => (x"50",x"c0",x"48",x"ef"),
   773 => (x"de",x"e4",x"c2",x"7e"),
   774 => (x"dc",x"c2",x"49",x"bf"),
   775 => (x"71",x"4a",x"bf",x"ce"),
   776 => (x"f7",x"fb",x"04",x"aa"),
   777 => (x"ff",x"e8",x"c2",x"87"),
   778 => (x"c8",x"c0",x"05",x"bf"),
   779 => (x"da",x"e4",x"c2",x"87"),
   780 => (x"f8",x"c1",x"02",x"bf"),
   781 => (x"ca",x"dc",x"c2",x"87"),
   782 => (x"df",x"ed",x"49",x"bf"),
   783 => (x"c2",x"49",x"70",x"87"),
   784 => (x"c4",x"59",x"ce",x"dc"),
   785 => (x"dc",x"c2",x"48",x"a6"),
   786 => (x"c2",x"78",x"bf",x"ca"),
   787 => (x"02",x"bf",x"da",x"e4"),
   788 => (x"c4",x"87",x"d8",x"c0"),
   789 => (x"ff",x"cf",x"49",x"66"),
   790 => (x"99",x"f8",x"ff",x"ff"),
   791 => (x"c5",x"c0",x"02",x"a9"),
   792 => (x"c0",x"4c",x"c0",x"87"),
   793 => (x"4c",x"c1",x"87",x"e1"),
   794 => (x"c4",x"87",x"dc",x"c0"),
   795 => (x"ff",x"cf",x"49",x"66"),
   796 => (x"02",x"a9",x"99",x"f8"),
   797 => (x"c8",x"87",x"c8",x"c0"),
   798 => (x"78",x"c0",x"48",x"a6"),
   799 => (x"c8",x"87",x"c5",x"c0"),
   800 => (x"78",x"c1",x"48",x"a6"),
   801 => (x"74",x"4c",x"66",x"c8"),
   802 => (x"e0",x"c0",x"05",x"9c"),
   803 => (x"49",x"66",x"c4",x"87"),
   804 => (x"e4",x"c2",x"89",x"c2"),
   805 => (x"91",x"4a",x"bf",x"d2"),
   806 => (x"bf",x"eb",x"e8",x"c2"),
   807 => (x"c6",x"dc",x"c2",x"4a"),
   808 => (x"78",x"a1",x"72",x"48"),
   809 => (x"48",x"ce",x"dc",x"c2"),
   810 => (x"df",x"f9",x"78",x"c0"),
   811 => (x"f4",x"48",x"c0",x"87"),
   812 => (x"87",x"e0",x"eb",x"8e"),
   813 => (x"00",x"00",x"00",x"00"),
   814 => (x"ff",x"ff",x"ff",x"ff"),
   815 => (x"00",x"00",x"0c",x"c4"),
   816 => (x"00",x"00",x"0c",x"cd"),
   817 => (x"33",x"54",x"41",x"46"),
   818 => (x"20",x"20",x"20",x"32"),
   819 => (x"54",x"41",x"46",x"00"),
   820 => (x"20",x"20",x"36",x"31"),
   821 => (x"ff",x"1e",x"00",x"20"),
   822 => (x"ff",x"c3",x"48",x"d4"),
   823 => (x"26",x"48",x"68",x"78"),
   824 => (x"d4",x"ff",x"1e",x"4f"),
   825 => (x"78",x"ff",x"c3",x"48"),
   826 => (x"c8",x"48",x"d0",x"ff"),
   827 => (x"d4",x"ff",x"78",x"e1"),
   828 => (x"c2",x"78",x"d4",x"48"),
   829 => (x"ff",x"48",x"c3",x"e9"),
   830 => (x"26",x"50",x"bf",x"d4"),
   831 => (x"d0",x"ff",x"1e",x"4f"),
   832 => (x"78",x"e0",x"c0",x"48"),
   833 => (x"ff",x"1e",x"4f",x"26"),
   834 => (x"49",x"70",x"87",x"cc"),
   835 => (x"87",x"c6",x"02",x"99"),
   836 => (x"05",x"a9",x"fb",x"c0"),
   837 => (x"48",x"71",x"87",x"f1"),
   838 => (x"5e",x"0e",x"4f",x"26"),
   839 => (x"71",x"0e",x"5c",x"5b"),
   840 => (x"fe",x"4c",x"c0",x"4b"),
   841 => (x"49",x"70",x"87",x"f0"),
   842 => (x"f9",x"c0",x"02",x"99"),
   843 => (x"a9",x"ec",x"c0",x"87"),
   844 => (x"87",x"f2",x"c0",x"02"),
   845 => (x"02",x"a9",x"fb",x"c0"),
   846 => (x"cc",x"87",x"eb",x"c0"),
   847 => (x"03",x"ac",x"b7",x"66"),
   848 => (x"66",x"d0",x"87",x"c7"),
   849 => (x"71",x"87",x"c2",x"02"),
   850 => (x"02",x"99",x"71",x"53"),
   851 => (x"84",x"c1",x"87",x"c2"),
   852 => (x"70",x"87",x"c3",x"fe"),
   853 => (x"cd",x"02",x"99",x"49"),
   854 => (x"a9",x"ec",x"c0",x"87"),
   855 => (x"c0",x"87",x"c7",x"02"),
   856 => (x"ff",x"05",x"a9",x"fb"),
   857 => (x"66",x"d0",x"87",x"d5"),
   858 => (x"c0",x"87",x"c3",x"02"),
   859 => (x"ec",x"c0",x"7b",x"97"),
   860 => (x"87",x"c4",x"05",x"a9"),
   861 => (x"87",x"c5",x"4a",x"74"),
   862 => (x"0a",x"c0",x"4a",x"74"),
   863 => (x"c2",x"48",x"72",x"8a"),
   864 => (x"26",x"4d",x"26",x"87"),
   865 => (x"26",x"4b",x"26",x"4c"),
   866 => (x"c9",x"fd",x"1e",x"4f"),
   867 => (x"c0",x"49",x"70",x"87"),
   868 => (x"04",x"a9",x"b7",x"f0"),
   869 => (x"f9",x"c0",x"87",x"ca"),
   870 => (x"c3",x"01",x"a9",x"b7"),
   871 => (x"89",x"f0",x"c0",x"87"),
   872 => (x"a9",x"b7",x"c1",x"c1"),
   873 => (x"c1",x"87",x"ca",x"04"),
   874 => (x"01",x"a9",x"b7",x"da"),
   875 => (x"f7",x"c0",x"87",x"c3"),
   876 => (x"26",x"48",x"71",x"89"),
   877 => (x"5b",x"5e",x"0e",x"4f"),
   878 => (x"4a",x"71",x"0e",x"5c"),
   879 => (x"72",x"4c",x"d4",x"ff"),
   880 => (x"87",x"ea",x"c0",x"49"),
   881 => (x"02",x"9b",x"4b",x"70"),
   882 => (x"8b",x"c1",x"87",x"c2"),
   883 => (x"c8",x"48",x"d0",x"ff"),
   884 => (x"d5",x"c1",x"78",x"c5"),
   885 => (x"c6",x"49",x"73",x"7c"),
   886 => (x"d1",x"e3",x"c1",x"31"),
   887 => (x"48",x"4a",x"bf",x"97"),
   888 => (x"7c",x"70",x"b0",x"71"),
   889 => (x"c4",x"48",x"d0",x"ff"),
   890 => (x"fe",x"48",x"73",x"78"),
   891 => (x"5e",x"0e",x"87",x"d5"),
   892 => (x"0e",x"5d",x"5c",x"5b"),
   893 => (x"4c",x"71",x"86",x"f8"),
   894 => (x"e4",x"fb",x"7e",x"c0"),
   895 => (x"c0",x"4b",x"c0",x"87"),
   896 => (x"bf",x"97",x"db",x"fa"),
   897 => (x"04",x"a9",x"c0",x"49"),
   898 => (x"f9",x"fb",x"87",x"cf"),
   899 => (x"c0",x"83",x"c1",x"87"),
   900 => (x"bf",x"97",x"db",x"fa"),
   901 => (x"f1",x"06",x"ab",x"49"),
   902 => (x"db",x"fa",x"c0",x"87"),
   903 => (x"cf",x"02",x"bf",x"97"),
   904 => (x"87",x"f2",x"fa",x"87"),
   905 => (x"02",x"99",x"49",x"70"),
   906 => (x"ec",x"c0",x"87",x"c6"),
   907 => (x"87",x"f1",x"05",x"a9"),
   908 => (x"e1",x"fa",x"4b",x"c0"),
   909 => (x"fa",x"4d",x"70",x"87"),
   910 => (x"a6",x"c8",x"87",x"dc"),
   911 => (x"87",x"d6",x"fa",x"58"),
   912 => (x"83",x"c1",x"4a",x"70"),
   913 => (x"97",x"49",x"a4",x"c8"),
   914 => (x"02",x"ad",x"49",x"69"),
   915 => (x"ff",x"c0",x"87",x"c7"),
   916 => (x"e7",x"c0",x"05",x"ad"),
   917 => (x"49",x"a4",x"c9",x"87"),
   918 => (x"c4",x"49",x"69",x"97"),
   919 => (x"c7",x"02",x"a9",x"66"),
   920 => (x"ff",x"c0",x"48",x"87"),
   921 => (x"87",x"d4",x"05",x"a8"),
   922 => (x"97",x"49",x"a4",x"ca"),
   923 => (x"02",x"aa",x"49",x"69"),
   924 => (x"ff",x"c0",x"87",x"c6"),
   925 => (x"87",x"c4",x"05",x"aa"),
   926 => (x"87",x"d0",x"7e",x"c1"),
   927 => (x"02",x"ad",x"ec",x"c0"),
   928 => (x"fb",x"c0",x"87",x"c6"),
   929 => (x"87",x"c4",x"05",x"ad"),
   930 => (x"7e",x"c1",x"4b",x"c0"),
   931 => (x"e1",x"fe",x"02",x"6e"),
   932 => (x"87",x"e9",x"f9",x"87"),
   933 => (x"8e",x"f8",x"48",x"73"),
   934 => (x"00",x"87",x"e6",x"fb"),
   935 => (x"5c",x"5b",x"5e",x"0e"),
   936 => (x"71",x"1e",x"0e",x"5d"),
   937 => (x"4b",x"d4",x"ff",x"4d"),
   938 => (x"e9",x"c2",x"1e",x"75"),
   939 => (x"fc",x"e6",x"49",x"c8"),
   940 => (x"70",x"86",x"c4",x"87"),
   941 => (x"d8",x"c3",x"02",x"98"),
   942 => (x"d0",x"e9",x"c2",x"87"),
   943 => (x"49",x"75",x"4c",x"bf"),
   944 => (x"ff",x"87",x"f2",x"fb"),
   945 => (x"c5",x"c8",x"48",x"d0"),
   946 => (x"7b",x"d6",x"c1",x"78"),
   947 => (x"a2",x"75",x"4a",x"c0"),
   948 => (x"c1",x"7b",x"11",x"49"),
   949 => (x"aa",x"b7",x"cb",x"82"),
   950 => (x"cc",x"87",x"f3",x"04"),
   951 => (x"7b",x"ff",x"c3",x"4a"),
   952 => (x"e0",x"c0",x"82",x"c1"),
   953 => (x"f4",x"04",x"aa",x"b7"),
   954 => (x"48",x"d0",x"ff",x"87"),
   955 => (x"ff",x"c3",x"78",x"c4"),
   956 => (x"78",x"c5",x"c8",x"7b"),
   957 => (x"c1",x"7b",x"d3",x"c1"),
   958 => (x"74",x"78",x"c4",x"7b"),
   959 => (x"ff",x"c1",x"02",x"9c"),
   960 => (x"d2",x"dc",x"c2",x"87"),
   961 => (x"4d",x"c0",x"c8",x"7e"),
   962 => (x"ac",x"b7",x"c0",x"8c"),
   963 => (x"c8",x"87",x"c6",x"03"),
   964 => (x"c0",x"4d",x"a4",x"c0"),
   965 => (x"ad",x"c0",x"c8",x"4c"),
   966 => (x"c2",x"87",x"dc",x"05"),
   967 => (x"bf",x"97",x"c3",x"e9"),
   968 => (x"02",x"99",x"d0",x"49"),
   969 => (x"1e",x"c0",x"87",x"d1"),
   970 => (x"49",x"c8",x"e9",x"c2"),
   971 => (x"c4",x"87",x"d3",x"e8"),
   972 => (x"4a",x"49",x"70",x"86"),
   973 => (x"c2",x"87",x"ee",x"c0"),
   974 => (x"c2",x"1e",x"d2",x"dc"),
   975 => (x"e8",x"49",x"c8",x"e9"),
   976 => (x"86",x"c4",x"87",x"c0"),
   977 => (x"ff",x"4a",x"49",x"70"),
   978 => (x"c5",x"c8",x"48",x"d0"),
   979 => (x"7b",x"d4",x"c1",x"78"),
   980 => (x"7b",x"bf",x"97",x"6e"),
   981 => (x"80",x"c1",x"48",x"6e"),
   982 => (x"8d",x"c1",x"7e",x"70"),
   983 => (x"87",x"f0",x"ff",x"05"),
   984 => (x"c4",x"48",x"d0",x"ff"),
   985 => (x"05",x"9a",x"72",x"78"),
   986 => (x"48",x"c0",x"87",x"c5"),
   987 => (x"c1",x"87",x"e4",x"c0"),
   988 => (x"c8",x"e9",x"c2",x"1e"),
   989 => (x"87",x"f0",x"e5",x"49"),
   990 => (x"9c",x"74",x"86",x"c4"),
   991 => (x"87",x"c1",x"fe",x"05"),
   992 => (x"c8",x"48",x"d0",x"ff"),
   993 => (x"d3",x"c1",x"78",x"c5"),
   994 => (x"c4",x"7b",x"c0",x"7b"),
   995 => (x"c2",x"48",x"c1",x"78"),
   996 => (x"26",x"48",x"c0",x"87"),
   997 => (x"4c",x"26",x"4d",x"26"),
   998 => (x"4f",x"26",x"4b",x"26"),
   999 => (x"5c",x"5b",x"5e",x"0e"),
  1000 => (x"71",x"1e",x"0e",x"5d"),
  1001 => (x"4d",x"4c",x"c0",x"4b"),
  1002 => (x"e8",x"c0",x"04",x"ab"),
  1003 => (x"ee",x"f7",x"c0",x"87"),
  1004 => (x"02",x"9d",x"75",x"1e"),
  1005 => (x"4a",x"c0",x"87",x"c4"),
  1006 => (x"4a",x"c1",x"87",x"c2"),
  1007 => (x"dc",x"ec",x"49",x"72"),
  1008 => (x"70",x"86",x"c4",x"87"),
  1009 => (x"6e",x"84",x"c1",x"7e"),
  1010 => (x"73",x"87",x"c2",x"05"),
  1011 => (x"73",x"85",x"c1",x"4c"),
  1012 => (x"d8",x"ff",x"06",x"ac"),
  1013 => (x"26",x"48",x"6e",x"87"),
  1014 => (x"0e",x"87",x"f9",x"fe"),
  1015 => (x"0e",x"5c",x"5b",x"5e"),
  1016 => (x"66",x"cc",x"4b",x"71"),
  1017 => (x"4c",x"87",x"d8",x"02"),
  1018 => (x"02",x"8c",x"f0",x"c0"),
  1019 => (x"4a",x"74",x"87",x"d8"),
  1020 => (x"d1",x"02",x"8a",x"c1"),
  1021 => (x"cd",x"02",x"8a",x"87"),
  1022 => (x"c9",x"02",x"8a",x"87"),
  1023 => (x"73",x"87",x"d9",x"87"),
  1024 => (x"87",x"d8",x"fa",x"49"),
  1025 => (x"1e",x"74",x"87",x"d2"),
  1026 => (x"d8",x"c1",x"49",x"c0"),
  1027 => (x"1e",x"74",x"87",x"cb"),
  1028 => (x"d8",x"c1",x"49",x"73"),
  1029 => (x"86",x"c8",x"87",x"c3"),
  1030 => (x"0e",x"87",x"fb",x"fd"),
  1031 => (x"5d",x"5c",x"5b",x"5e"),
  1032 => (x"4c",x"71",x"1e",x"0e"),
  1033 => (x"c2",x"91",x"de",x"49"),
  1034 => (x"71",x"4d",x"f0",x"e9"),
  1035 => (x"02",x"6d",x"97",x"85"),
  1036 => (x"c2",x"87",x"dc",x"c1"),
  1037 => (x"4a",x"bf",x"dc",x"e9"),
  1038 => (x"49",x"72",x"82",x"74"),
  1039 => (x"70",x"87",x"dd",x"fd"),
  1040 => (x"c0",x"02",x"6e",x"7e"),
  1041 => (x"e9",x"c2",x"87",x"f2"),
  1042 => (x"4a",x"6e",x"4b",x"e4"),
  1043 => (x"c1",x"ff",x"49",x"cb"),
  1044 => (x"4b",x"74",x"87",x"d6"),
  1045 => (x"e3",x"c1",x"93",x"cb"),
  1046 => (x"83",x"c4",x"83",x"e1"),
  1047 => (x"7b",x"d3",x"c2",x"c1"),
  1048 => (x"c2",x"c1",x"49",x"74"),
  1049 => (x"7b",x"75",x"87",x"cd"),
  1050 => (x"97",x"d2",x"e3",x"c1"),
  1051 => (x"c2",x"1e",x"49",x"bf"),
  1052 => (x"fd",x"49",x"e4",x"e9"),
  1053 => (x"86",x"c4",x"87",x"e5"),
  1054 => (x"c1",x"c1",x"49",x"74"),
  1055 => (x"49",x"c0",x"87",x"f5"),
  1056 => (x"87",x"d4",x"c3",x"c1"),
  1057 => (x"48",x"c4",x"e9",x"c2"),
  1058 => (x"49",x"c1",x"78",x"c0"),
  1059 => (x"26",x"87",x"c1",x"dd"),
  1060 => (x"4c",x"87",x"c1",x"fc"),
  1061 => (x"69",x"64",x"61",x"6f"),
  1062 => (x"2e",x"2e",x"67",x"6e"),
  1063 => (x"5e",x"0e",x"00",x"2e"),
  1064 => (x"71",x"0e",x"5c",x"5b"),
  1065 => (x"e9",x"c2",x"4a",x"4b"),
  1066 => (x"72",x"82",x"bf",x"dc"),
  1067 => (x"87",x"ec",x"fb",x"49"),
  1068 => (x"02",x"9c",x"4c",x"70"),
  1069 => (x"e7",x"49",x"87",x"c4"),
  1070 => (x"e9",x"c2",x"87",x"eb"),
  1071 => (x"78",x"c0",x"48",x"dc"),
  1072 => (x"cb",x"dc",x"49",x"c1"),
  1073 => (x"87",x"ce",x"fb",x"87"),
  1074 => (x"5c",x"5b",x"5e",x"0e"),
  1075 => (x"86",x"f4",x"0e",x"5d"),
  1076 => (x"4d",x"d2",x"dc",x"c2"),
  1077 => (x"a6",x"c4",x"4c",x"c0"),
  1078 => (x"c2",x"78",x"c0",x"48"),
  1079 => (x"49",x"bf",x"dc",x"e9"),
  1080 => (x"c1",x"06",x"a9",x"c0"),
  1081 => (x"dc",x"c2",x"87",x"c1"),
  1082 => (x"02",x"98",x"48",x"d2"),
  1083 => (x"c0",x"87",x"f8",x"c0"),
  1084 => (x"c8",x"1e",x"ee",x"f7"),
  1085 => (x"87",x"c7",x"02",x"66"),
  1086 => (x"c0",x"48",x"a6",x"c4"),
  1087 => (x"c4",x"87",x"c5",x"78"),
  1088 => (x"78",x"c1",x"48",x"a6"),
  1089 => (x"e7",x"49",x"66",x"c4"),
  1090 => (x"86",x"c4",x"87",x"d3"),
  1091 => (x"84",x"c1",x"4d",x"70"),
  1092 => (x"c1",x"48",x"66",x"c4"),
  1093 => (x"58",x"a6",x"c8",x"80"),
  1094 => (x"bf",x"dc",x"e9",x"c2"),
  1095 => (x"c6",x"03",x"ac",x"49"),
  1096 => (x"05",x"9d",x"75",x"87"),
  1097 => (x"c0",x"87",x"c8",x"ff"),
  1098 => (x"02",x"9d",x"75",x"4c"),
  1099 => (x"c0",x"87",x"e0",x"c3"),
  1100 => (x"c8",x"1e",x"ee",x"f7"),
  1101 => (x"87",x"c7",x"02",x"66"),
  1102 => (x"c0",x"48",x"a6",x"cc"),
  1103 => (x"cc",x"87",x"c5",x"78"),
  1104 => (x"78",x"c1",x"48",x"a6"),
  1105 => (x"e6",x"49",x"66",x"cc"),
  1106 => (x"86",x"c4",x"87",x"d3"),
  1107 => (x"02",x"6e",x"7e",x"70"),
  1108 => (x"6e",x"87",x"e9",x"c2"),
  1109 => (x"97",x"81",x"cb",x"49"),
  1110 => (x"99",x"d0",x"49",x"69"),
  1111 => (x"87",x"d6",x"c1",x"02"),
  1112 => (x"4a",x"de",x"c2",x"c1"),
  1113 => (x"91",x"cb",x"49",x"74"),
  1114 => (x"81",x"e1",x"e3",x"c1"),
  1115 => (x"81",x"c8",x"79",x"72"),
  1116 => (x"74",x"51",x"ff",x"c3"),
  1117 => (x"c2",x"91",x"de",x"49"),
  1118 => (x"71",x"4d",x"f0",x"e9"),
  1119 => (x"97",x"c1",x"c2",x"85"),
  1120 => (x"49",x"a5",x"c1",x"7d"),
  1121 => (x"c2",x"51",x"e0",x"c0"),
  1122 => (x"bf",x"97",x"e2",x"e4"),
  1123 => (x"c1",x"87",x"d2",x"02"),
  1124 => (x"4b",x"a5",x"c2",x"84"),
  1125 => (x"4a",x"e2",x"e4",x"c2"),
  1126 => (x"fc",x"fe",x"49",x"db"),
  1127 => (x"db",x"c1",x"87",x"ca"),
  1128 => (x"49",x"a5",x"cd",x"87"),
  1129 => (x"84",x"c1",x"51",x"c0"),
  1130 => (x"6e",x"4b",x"a5",x"c2"),
  1131 => (x"fe",x"49",x"cb",x"4a"),
  1132 => (x"c1",x"87",x"f5",x"fb"),
  1133 => (x"c0",x"c1",x"87",x"c6"),
  1134 => (x"49",x"74",x"4a",x"db"),
  1135 => (x"e3",x"c1",x"91",x"cb"),
  1136 => (x"79",x"72",x"81",x"e1"),
  1137 => (x"97",x"e2",x"e4",x"c2"),
  1138 => (x"87",x"d8",x"02",x"bf"),
  1139 => (x"91",x"de",x"49",x"74"),
  1140 => (x"e9",x"c2",x"84",x"c1"),
  1141 => (x"83",x"71",x"4b",x"f0"),
  1142 => (x"4a",x"e2",x"e4",x"c2"),
  1143 => (x"fb",x"fe",x"49",x"dd"),
  1144 => (x"87",x"d8",x"87",x"c6"),
  1145 => (x"93",x"de",x"4b",x"74"),
  1146 => (x"83",x"f0",x"e9",x"c2"),
  1147 => (x"c0",x"49",x"a3",x"cb"),
  1148 => (x"73",x"84",x"c1",x"51"),
  1149 => (x"49",x"cb",x"4a",x"6e"),
  1150 => (x"87",x"ec",x"fa",x"fe"),
  1151 => (x"c1",x"48",x"66",x"c4"),
  1152 => (x"58",x"a6",x"c8",x"80"),
  1153 => (x"c0",x"03",x"ac",x"c7"),
  1154 => (x"05",x"6e",x"87",x"c5"),
  1155 => (x"74",x"87",x"e0",x"fc"),
  1156 => (x"f5",x"8e",x"f4",x"48"),
  1157 => (x"73",x"1e",x"87",x"fe"),
  1158 => (x"49",x"4b",x"71",x"1e"),
  1159 => (x"e3",x"c1",x"91",x"cb"),
  1160 => (x"a1",x"c8",x"81",x"e1"),
  1161 => (x"d1",x"e3",x"c1",x"4a"),
  1162 => (x"c9",x"50",x"12",x"48"),
  1163 => (x"fa",x"c0",x"4a",x"a1"),
  1164 => (x"50",x"12",x"48",x"db"),
  1165 => (x"e3",x"c1",x"81",x"ca"),
  1166 => (x"50",x"11",x"48",x"d2"),
  1167 => (x"97",x"d2",x"e3",x"c1"),
  1168 => (x"c0",x"1e",x"49",x"bf"),
  1169 => (x"87",x"d3",x"f6",x"49"),
  1170 => (x"48",x"c4",x"e9",x"c2"),
  1171 => (x"49",x"c1",x"78",x"de"),
  1172 => (x"26",x"87",x"fd",x"d5"),
  1173 => (x"1e",x"87",x"c1",x"f5"),
  1174 => (x"cb",x"49",x"4a",x"71"),
  1175 => (x"e1",x"e3",x"c1",x"91"),
  1176 => (x"11",x"81",x"c8",x"81"),
  1177 => (x"c8",x"e9",x"c2",x"48"),
  1178 => (x"dc",x"e9",x"c2",x"58"),
  1179 => (x"c1",x"78",x"c0",x"48"),
  1180 => (x"87",x"dc",x"d5",x"49"),
  1181 => (x"c0",x"1e",x"4f",x"26"),
  1182 => (x"db",x"fb",x"c0",x"49"),
  1183 => (x"1e",x"4f",x"26",x"87"),
  1184 => (x"d2",x"02",x"99",x"71"),
  1185 => (x"f6",x"e4",x"c1",x"87"),
  1186 => (x"f7",x"50",x"c0",x"48"),
  1187 => (x"d7",x"c9",x"c1",x"80"),
  1188 => (x"da",x"e3",x"c1",x"40"),
  1189 => (x"c1",x"87",x"ce",x"78"),
  1190 => (x"c1",x"48",x"f2",x"e4"),
  1191 => (x"fc",x"78",x"d3",x"e3"),
  1192 => (x"f6",x"c9",x"c1",x"80"),
  1193 => (x"0e",x"4f",x"26",x"78"),
  1194 => (x"0e",x"5c",x"5b",x"5e"),
  1195 => (x"cb",x"4a",x"4c",x"71"),
  1196 => (x"e1",x"e3",x"c1",x"92"),
  1197 => (x"49",x"a2",x"c8",x"82"),
  1198 => (x"97",x"4b",x"a2",x"c9"),
  1199 => (x"97",x"1e",x"4b",x"6b"),
  1200 => (x"ca",x"1e",x"49",x"69"),
  1201 => (x"c0",x"49",x"12",x"82"),
  1202 => (x"c0",x"87",x"d6",x"e6"),
  1203 => (x"87",x"c0",x"d4",x"49"),
  1204 => (x"f8",x"c0",x"49",x"74"),
  1205 => (x"8e",x"f8",x"87",x"dd"),
  1206 => (x"1e",x"87",x"fb",x"f2"),
  1207 => (x"4b",x"71",x"1e",x"73"),
  1208 => (x"87",x"c3",x"ff",x"49"),
  1209 => (x"fe",x"fe",x"49",x"73"),
  1210 => (x"87",x"ec",x"f2",x"87"),
  1211 => (x"71",x"1e",x"73",x"1e"),
  1212 => (x"4a",x"a3",x"c6",x"4b"),
  1213 => (x"c1",x"87",x"db",x"02"),
  1214 => (x"87",x"d6",x"02",x"8a"),
  1215 => (x"da",x"c1",x"02",x"8a"),
  1216 => (x"c0",x"02",x"8a",x"87"),
  1217 => (x"02",x"8a",x"87",x"fc"),
  1218 => (x"8a",x"87",x"e1",x"c0"),
  1219 => (x"c1",x"87",x"cb",x"02"),
  1220 => (x"49",x"c7",x"87",x"db"),
  1221 => (x"c1",x"87",x"c0",x"fd"),
  1222 => (x"e9",x"c2",x"87",x"de"),
  1223 => (x"c1",x"02",x"bf",x"dc"),
  1224 => (x"c1",x"48",x"87",x"cb"),
  1225 => (x"e0",x"e9",x"c2",x"88"),
  1226 => (x"87",x"c1",x"c1",x"58"),
  1227 => (x"bf",x"e0",x"e9",x"c2"),
  1228 => (x"87",x"f9",x"c0",x"02"),
  1229 => (x"bf",x"dc",x"e9",x"c2"),
  1230 => (x"c2",x"80",x"c1",x"48"),
  1231 => (x"c0",x"58",x"e0",x"e9"),
  1232 => (x"e9",x"c2",x"87",x"eb"),
  1233 => (x"c6",x"49",x"bf",x"dc"),
  1234 => (x"e0",x"e9",x"c2",x"89"),
  1235 => (x"a9",x"b7",x"c0",x"59"),
  1236 => (x"c2",x"87",x"da",x"03"),
  1237 => (x"c0",x"48",x"dc",x"e9"),
  1238 => (x"c2",x"87",x"d2",x"78"),
  1239 => (x"02",x"bf",x"e0",x"e9"),
  1240 => (x"e9",x"c2",x"87",x"cb"),
  1241 => (x"c6",x"48",x"bf",x"dc"),
  1242 => (x"e0",x"e9",x"c2",x"80"),
  1243 => (x"d1",x"49",x"c0",x"58"),
  1244 => (x"49",x"73",x"87",x"de"),
  1245 => (x"87",x"fb",x"f5",x"c0"),
  1246 => (x"0e",x"87",x"dd",x"f0"),
  1247 => (x"0e",x"5c",x"5b",x"5e"),
  1248 => (x"66",x"cc",x"4c",x"71"),
  1249 => (x"cb",x"4b",x"74",x"1e"),
  1250 => (x"e1",x"e3",x"c1",x"93"),
  1251 => (x"4a",x"a3",x"c4",x"83"),
  1252 => (x"f4",x"fe",x"49",x"6a"),
  1253 => (x"c8",x"c1",x"87",x"e2"),
  1254 => (x"a3",x"c8",x"7b",x"d6"),
  1255 => (x"51",x"66",x"d4",x"49"),
  1256 => (x"d8",x"49",x"a3",x"c9"),
  1257 => (x"a3",x"ca",x"51",x"66"),
  1258 => (x"51",x"66",x"dc",x"49"),
  1259 => (x"87",x"e6",x"ef",x"26"),
  1260 => (x"5c",x"5b",x"5e",x"0e"),
  1261 => (x"d0",x"ff",x"0e",x"5d"),
  1262 => (x"59",x"a6",x"d8",x"86"),
  1263 => (x"c0",x"48",x"a6",x"c4"),
  1264 => (x"c1",x"80",x"c4",x"78"),
  1265 => (x"c4",x"78",x"66",x"c4"),
  1266 => (x"c4",x"78",x"c1",x"80"),
  1267 => (x"c2",x"78",x"c1",x"80"),
  1268 => (x"c1",x"48",x"e0",x"e9"),
  1269 => (x"c4",x"e9",x"c2",x"78"),
  1270 => (x"a8",x"de",x"48",x"bf"),
  1271 => (x"f3",x"87",x"cb",x"05"),
  1272 => (x"49",x"70",x"87",x"e6"),
  1273 => (x"ce",x"59",x"a6",x"c8"),
  1274 => (x"f4",x"e3",x"87",x"ee"),
  1275 => (x"87",x"d6",x"e4",x"87"),
  1276 => (x"70",x"87",x"e3",x"e3"),
  1277 => (x"ac",x"fb",x"c0",x"4c"),
  1278 => (x"87",x"d0",x"c1",x"02"),
  1279 => (x"c1",x"05",x"66",x"d4"),
  1280 => (x"1e",x"c0",x"87",x"c2"),
  1281 => (x"c1",x"1e",x"c1",x"1e"),
  1282 => (x"c0",x"1e",x"d4",x"e5"),
  1283 => (x"87",x"eb",x"fd",x"49"),
  1284 => (x"4a",x"66",x"d0",x"c1"),
  1285 => (x"49",x"6a",x"82",x"c4"),
  1286 => (x"51",x"74",x"81",x"c7"),
  1287 => (x"1e",x"d8",x"1e",x"c1"),
  1288 => (x"81",x"c8",x"49",x"6a"),
  1289 => (x"d8",x"87",x"f3",x"e3"),
  1290 => (x"66",x"c4",x"c1",x"86"),
  1291 => (x"01",x"a8",x"c0",x"48"),
  1292 => (x"a6",x"c4",x"87",x"c7"),
  1293 => (x"ce",x"78",x"c1",x"48"),
  1294 => (x"66",x"c4",x"c1",x"87"),
  1295 => (x"cc",x"88",x"c1",x"48"),
  1296 => (x"87",x"c3",x"58",x"a6"),
  1297 => (x"cc",x"87",x"ff",x"e2"),
  1298 => (x"78",x"c2",x"48",x"a6"),
  1299 => (x"cd",x"02",x"9c",x"74"),
  1300 => (x"66",x"c4",x"87",x"c2"),
  1301 => (x"66",x"c8",x"c1",x"48"),
  1302 => (x"f7",x"cc",x"03",x"a8"),
  1303 => (x"48",x"a6",x"d8",x"87"),
  1304 => (x"80",x"c4",x"78",x"c0"),
  1305 => (x"ed",x"e1",x"78",x"c0"),
  1306 => (x"c1",x"4c",x"70",x"87"),
  1307 => (x"c2",x"05",x"ac",x"d0"),
  1308 => (x"66",x"dc",x"87",x"d8"),
  1309 => (x"87",x"d1",x"e4",x"7e"),
  1310 => (x"e0",x"c0",x"49",x"70"),
  1311 => (x"d5",x"e1",x"59",x"a6"),
  1312 => (x"c0",x"4c",x"70",x"87"),
  1313 => (x"c1",x"05",x"ac",x"ec"),
  1314 => (x"66",x"c4",x"87",x"eb"),
  1315 => (x"c1",x"91",x"cb",x"49"),
  1316 => (x"c4",x"81",x"66",x"c0"),
  1317 => (x"4d",x"6a",x"4a",x"a1"),
  1318 => (x"dc",x"4a",x"a1",x"c8"),
  1319 => (x"c9",x"c1",x"52",x"66"),
  1320 => (x"f1",x"e0",x"79",x"d7"),
  1321 => (x"9c",x"4c",x"70",x"87"),
  1322 => (x"c0",x"87",x"d8",x"02"),
  1323 => (x"d2",x"02",x"ac",x"fb"),
  1324 => (x"e0",x"55",x"74",x"87"),
  1325 => (x"4c",x"70",x"87",x"e0"),
  1326 => (x"87",x"c7",x"02",x"9c"),
  1327 => (x"05",x"ac",x"fb",x"c0"),
  1328 => (x"c0",x"87",x"ee",x"ff"),
  1329 => (x"c1",x"c2",x"55",x"e0"),
  1330 => (x"7d",x"97",x"c0",x"55"),
  1331 => (x"6e",x"49",x"66",x"d4"),
  1332 => (x"87",x"db",x"05",x"a9"),
  1333 => (x"c8",x"48",x"66",x"c4"),
  1334 => (x"ca",x"04",x"a8",x"66"),
  1335 => (x"48",x"66",x"c4",x"87"),
  1336 => (x"a6",x"c8",x"80",x"c1"),
  1337 => (x"c8",x"87",x"c8",x"58"),
  1338 => (x"88",x"c1",x"48",x"66"),
  1339 => (x"ff",x"58",x"a6",x"cc"),
  1340 => (x"70",x"87",x"e3",x"df"),
  1341 => (x"ac",x"d0",x"c1",x"4c"),
  1342 => (x"d0",x"87",x"c8",x"05"),
  1343 => (x"80",x"c1",x"48",x"66"),
  1344 => (x"c1",x"58",x"a6",x"d4"),
  1345 => (x"fd",x"02",x"ac",x"d0"),
  1346 => (x"e0",x"c0",x"87",x"e8"),
  1347 => (x"66",x"d4",x"48",x"a6"),
  1348 => (x"48",x"66",x"dc",x"78"),
  1349 => (x"a8",x"66",x"e0",x"c0"),
  1350 => (x"87",x"ca",x"c9",x"05"),
  1351 => (x"48",x"a6",x"e4",x"c0"),
  1352 => (x"74",x"7e",x"78",x"c0"),
  1353 => (x"88",x"fb",x"c0",x"48"),
  1354 => (x"58",x"a6",x"ec",x"c0"),
  1355 => (x"c8",x"02",x"98",x"70"),
  1356 => (x"cb",x"48",x"87",x"cf"),
  1357 => (x"a6",x"ec",x"c0",x"88"),
  1358 => (x"02",x"98",x"70",x"58"),
  1359 => (x"48",x"87",x"d2",x"c1"),
  1360 => (x"ec",x"c0",x"88",x"c9"),
  1361 => (x"98",x"70",x"58",x"a6"),
  1362 => (x"87",x"db",x"c3",x"02"),
  1363 => (x"c0",x"88",x"c4",x"48"),
  1364 => (x"70",x"58",x"a6",x"ec"),
  1365 => (x"87",x"d0",x"02",x"98"),
  1366 => (x"c0",x"88",x"c1",x"48"),
  1367 => (x"70",x"58",x"a6",x"ec"),
  1368 => (x"c2",x"c3",x"02",x"98"),
  1369 => (x"87",x"d3",x"c7",x"87"),
  1370 => (x"c0",x"48",x"a6",x"d8"),
  1371 => (x"dd",x"ff",x"78",x"f0"),
  1372 => (x"4c",x"70",x"87",x"e4"),
  1373 => (x"02",x"ac",x"ec",x"c0"),
  1374 => (x"dc",x"87",x"c3",x"c0"),
  1375 => (x"ec",x"c0",x"5c",x"a6"),
  1376 => (x"87",x"cd",x"02",x"ac"),
  1377 => (x"87",x"ce",x"dd",x"ff"),
  1378 => (x"ec",x"c0",x"4c",x"70"),
  1379 => (x"f3",x"ff",x"05",x"ac"),
  1380 => (x"ac",x"ec",x"c0",x"87"),
  1381 => (x"87",x"c4",x"c0",x"02"),
  1382 => (x"87",x"fa",x"dc",x"ff"),
  1383 => (x"d4",x"1e",x"66",x"d8"),
  1384 => (x"d4",x"1e",x"49",x"66"),
  1385 => (x"c1",x"1e",x"49",x"66"),
  1386 => (x"d4",x"1e",x"d4",x"e5"),
  1387 => (x"ca",x"f7",x"49",x"66"),
  1388 => (x"ca",x"1e",x"c0",x"87"),
  1389 => (x"49",x"66",x"dc",x"1e"),
  1390 => (x"d8",x"c1",x"91",x"cb"),
  1391 => (x"a6",x"d8",x"81",x"66"),
  1392 => (x"78",x"a1",x"c4",x"48"),
  1393 => (x"49",x"bf",x"66",x"d8"),
  1394 => (x"87",x"ce",x"dd",x"ff"),
  1395 => (x"b7",x"c0",x"86",x"d8"),
  1396 => (x"c5",x"c1",x"06",x"a8"),
  1397 => (x"de",x"1e",x"c1",x"87"),
  1398 => (x"bf",x"66",x"c8",x"1e"),
  1399 => (x"f9",x"dc",x"ff",x"49"),
  1400 => (x"70",x"86",x"c8",x"87"),
  1401 => (x"08",x"c0",x"48",x"49"),
  1402 => (x"58",x"a6",x"dc",x"88"),
  1403 => (x"06",x"a8",x"b7",x"c0"),
  1404 => (x"d8",x"87",x"e7",x"c0"),
  1405 => (x"b7",x"dd",x"48",x"66"),
  1406 => (x"87",x"de",x"03",x"a8"),
  1407 => (x"d8",x"49",x"bf",x"6e"),
  1408 => (x"e0",x"c0",x"81",x"66"),
  1409 => (x"49",x"66",x"d8",x"51"),
  1410 => (x"bf",x"6e",x"81",x"c1"),
  1411 => (x"51",x"c1",x"c2",x"81"),
  1412 => (x"c2",x"49",x"66",x"d8"),
  1413 => (x"81",x"bf",x"6e",x"81"),
  1414 => (x"66",x"cc",x"51",x"c0"),
  1415 => (x"d0",x"80",x"c1",x"48"),
  1416 => (x"7e",x"c1",x"58",x"a6"),
  1417 => (x"ff",x"87",x"da",x"c4"),
  1418 => (x"dc",x"87",x"de",x"dd"),
  1419 => (x"dd",x"ff",x"58",x"a6"),
  1420 => (x"ec",x"c0",x"87",x"d7"),
  1421 => (x"ec",x"c0",x"58",x"a6"),
  1422 => (x"ca",x"c0",x"05",x"a8"),
  1423 => (x"a6",x"e8",x"c0",x"87"),
  1424 => (x"78",x"66",x"d8",x"48"),
  1425 => (x"ff",x"87",x"c4",x"c0"),
  1426 => (x"c4",x"87",x"cb",x"da"),
  1427 => (x"91",x"cb",x"49",x"66"),
  1428 => (x"48",x"66",x"c0",x"c1"),
  1429 => (x"7e",x"70",x"80",x"71"),
  1430 => (x"82",x"c8",x"4a",x"6e"),
  1431 => (x"81",x"ca",x"49",x"6e"),
  1432 => (x"c0",x"51",x"66",x"d8"),
  1433 => (x"c1",x"49",x"66",x"e8"),
  1434 => (x"89",x"66",x"d8",x"81"),
  1435 => (x"30",x"71",x"48",x"c1"),
  1436 => (x"89",x"c1",x"49",x"70"),
  1437 => (x"c2",x"7a",x"97",x"71"),
  1438 => (x"49",x"bf",x"cc",x"ed"),
  1439 => (x"97",x"29",x"66",x"d8"),
  1440 => (x"71",x"48",x"4a",x"6a"),
  1441 => (x"a6",x"f0",x"c0",x"98"),
  1442 => (x"c4",x"49",x"6e",x"58"),
  1443 => (x"c0",x"4d",x"69",x"81"),
  1444 => (x"dc",x"48",x"66",x"e0"),
  1445 => (x"c0",x"02",x"a8",x"66"),
  1446 => (x"a6",x"d8",x"87",x"c8"),
  1447 => (x"c0",x"78",x"c0",x"48"),
  1448 => (x"a6",x"d8",x"87",x"c5"),
  1449 => (x"d8",x"78",x"c1",x"48"),
  1450 => (x"e0",x"c0",x"1e",x"66"),
  1451 => (x"ff",x"49",x"75",x"1e"),
  1452 => (x"c8",x"87",x"e7",x"d9"),
  1453 => (x"c0",x"4c",x"70",x"86"),
  1454 => (x"c1",x"06",x"ac",x"b7"),
  1455 => (x"85",x"74",x"87",x"d4"),
  1456 => (x"74",x"49",x"e0",x"c0"),
  1457 => (x"c1",x"4b",x"75",x"89"),
  1458 => (x"71",x"4a",x"cd",x"df"),
  1459 => (x"87",x"d8",x"e7",x"fe"),
  1460 => (x"e4",x"c0",x"85",x"c2"),
  1461 => (x"80",x"c1",x"48",x"66"),
  1462 => (x"58",x"a6",x"e8",x"c0"),
  1463 => (x"49",x"66",x"ec",x"c0"),
  1464 => (x"a9",x"70",x"81",x"c1"),
  1465 => (x"87",x"c8",x"c0",x"02"),
  1466 => (x"c0",x"48",x"a6",x"d8"),
  1467 => (x"87",x"c5",x"c0",x"78"),
  1468 => (x"c1",x"48",x"a6",x"d8"),
  1469 => (x"1e",x"66",x"d8",x"78"),
  1470 => (x"c0",x"49",x"a4",x"c2"),
  1471 => (x"88",x"71",x"48",x"e0"),
  1472 => (x"75",x"1e",x"49",x"70"),
  1473 => (x"d1",x"d8",x"ff",x"49"),
  1474 => (x"c0",x"86",x"c8",x"87"),
  1475 => (x"ff",x"01",x"a8",x"b7"),
  1476 => (x"e4",x"c0",x"87",x"c0"),
  1477 => (x"d1",x"c0",x"02",x"66"),
  1478 => (x"c9",x"49",x"6e",x"87"),
  1479 => (x"66",x"e4",x"c0",x"81"),
  1480 => (x"c1",x"48",x"6e",x"51"),
  1481 => (x"c0",x"78",x"e7",x"ca"),
  1482 => (x"49",x"6e",x"87",x"cc"),
  1483 => (x"51",x"c2",x"81",x"c9"),
  1484 => (x"cb",x"c1",x"48",x"6e"),
  1485 => (x"7e",x"c1",x"78",x"db"),
  1486 => (x"ff",x"87",x"c6",x"c0"),
  1487 => (x"70",x"87",x"c7",x"d7"),
  1488 => (x"c0",x"02",x"6e",x"4c"),
  1489 => (x"66",x"c4",x"87",x"f5"),
  1490 => (x"a8",x"66",x"c8",x"48"),
  1491 => (x"87",x"cb",x"c0",x"04"),
  1492 => (x"c1",x"48",x"66",x"c4"),
  1493 => (x"58",x"a6",x"c8",x"80"),
  1494 => (x"c8",x"87",x"e0",x"c0"),
  1495 => (x"88",x"c1",x"48",x"66"),
  1496 => (x"c0",x"58",x"a6",x"cc"),
  1497 => (x"c6",x"c1",x"87",x"d5"),
  1498 => (x"c8",x"c0",x"05",x"ac"),
  1499 => (x"48",x"66",x"cc",x"87"),
  1500 => (x"a6",x"d0",x"80",x"c1"),
  1501 => (x"cd",x"d6",x"ff",x"58"),
  1502 => (x"d0",x"4c",x"70",x"87"),
  1503 => (x"80",x"c1",x"48",x"66"),
  1504 => (x"74",x"58",x"a6",x"d4"),
  1505 => (x"cb",x"c0",x"02",x"9c"),
  1506 => (x"48",x"66",x"c4",x"87"),
  1507 => (x"a8",x"66",x"c8",x"c1"),
  1508 => (x"87",x"c9",x"f3",x"04"),
  1509 => (x"87",x"e5",x"d5",x"ff"),
  1510 => (x"c7",x"48",x"66",x"c4"),
  1511 => (x"e5",x"c0",x"03",x"a8"),
  1512 => (x"e0",x"e9",x"c2",x"87"),
  1513 => (x"c4",x"78",x"c0",x"48"),
  1514 => (x"91",x"cb",x"49",x"66"),
  1515 => (x"81",x"66",x"c0",x"c1"),
  1516 => (x"6a",x"4a",x"a1",x"c4"),
  1517 => (x"79",x"52",x"c0",x"4a"),
  1518 => (x"c1",x"48",x"66",x"c4"),
  1519 => (x"58",x"a6",x"c8",x"80"),
  1520 => (x"ff",x"04",x"a8",x"c7"),
  1521 => (x"d0",x"ff",x"87",x"db"),
  1522 => (x"c7",x"df",x"ff",x"8e"),
  1523 => (x"00",x"20",x"3a",x"87"),
  1524 => (x"71",x"1e",x"73",x"1e"),
  1525 => (x"c6",x"02",x"9b",x"4b"),
  1526 => (x"dc",x"e9",x"c2",x"87"),
  1527 => (x"c7",x"78",x"c0",x"48"),
  1528 => (x"dc",x"e9",x"c2",x"1e"),
  1529 => (x"c1",x"1e",x"49",x"bf"),
  1530 => (x"c2",x"1e",x"e1",x"e3"),
  1531 => (x"49",x"bf",x"c4",x"e9"),
  1532 => (x"cc",x"87",x"fd",x"ee"),
  1533 => (x"c4",x"e9",x"c2",x"86"),
  1534 => (x"c2",x"ea",x"49",x"bf"),
  1535 => (x"02",x"9b",x"73",x"87"),
  1536 => (x"e3",x"c1",x"87",x"c8"),
  1537 => (x"e4",x"c0",x"49",x"e1"),
  1538 => (x"de",x"ff",x"87",x"fb"),
  1539 => (x"73",x"1e",x"87",x"ca"),
  1540 => (x"c1",x"4b",x"c0",x"1e"),
  1541 => (x"c0",x"48",x"d1",x"e3"),
  1542 => (x"c4",x"e5",x"c1",x"50"),
  1543 => (x"d9",x"ff",x"49",x"bf"),
  1544 => (x"98",x"70",x"87",x"fa"),
  1545 => (x"c1",x"87",x"c4",x"05"),
  1546 => (x"73",x"4b",x"f1",x"e0"),
  1547 => (x"e7",x"dd",x"ff",x"48"),
  1548 => (x"4d",x"4f",x"52",x"87"),
  1549 => (x"61",x"6f",x"6c",x"20"),
  1550 => (x"67",x"6e",x"69",x"64"),
  1551 => (x"69",x"61",x"66",x"20"),
  1552 => (x"00",x"64",x"65",x"6c"),
  1553 => (x"87",x"eb",x"c7",x"1e"),
  1554 => (x"c3",x"fe",x"49",x"c1"),
  1555 => (x"cc",x"ea",x"fe",x"87"),
  1556 => (x"02",x"98",x"70",x"87"),
  1557 => (x"f3",x"fe",x"87",x"cd"),
  1558 => (x"98",x"70",x"87",x"c7"),
  1559 => (x"c1",x"87",x"c4",x"02"),
  1560 => (x"c0",x"87",x"c2",x"4a"),
  1561 => (x"05",x"9a",x"72",x"4a"),
  1562 => (x"1e",x"c0",x"87",x"ce"),
  1563 => (x"49",x"d8",x"e2",x"c1"),
  1564 => (x"87",x"df",x"ef",x"c0"),
  1565 => (x"87",x"fe",x"86",x"c4"),
  1566 => (x"87",x"c7",x"f9",x"c0"),
  1567 => (x"e2",x"c1",x"1e",x"c0"),
  1568 => (x"ef",x"c0",x"49",x"e3"),
  1569 => (x"1e",x"c0",x"87",x"cd"),
  1570 => (x"70",x"87",x"c3",x"fe"),
  1571 => (x"c2",x"ef",x"c0",x"49"),
  1572 => (x"87",x"de",x"c3",x"87"),
  1573 => (x"4f",x"26",x"8e",x"f8"),
  1574 => (x"66",x"20",x"44",x"53"),
  1575 => (x"65",x"6c",x"69",x"61"),
  1576 => (x"42",x"00",x"2e",x"64"),
  1577 => (x"69",x"74",x"6f",x"6f"),
  1578 => (x"2e",x"2e",x"67",x"6e"),
  1579 => (x"c0",x"1e",x"00",x"2e"),
  1580 => (x"c0",x"87",x"ee",x"e6"),
  1581 => (x"f6",x"87",x"d2",x"f2"),
  1582 => (x"1e",x"4f",x"26",x"87"),
  1583 => (x"48",x"dc",x"e9",x"c2"),
  1584 => (x"e9",x"c2",x"78",x"c0"),
  1585 => (x"78",x"c0",x"48",x"c4"),
  1586 => (x"e1",x"87",x"f9",x"fd"),
  1587 => (x"26",x"48",x"c0",x"87"),
  1588 => (x"80",x"00",x"00",x"4f"),
  1589 => (x"69",x"78",x"45",x"20"),
  1590 => (x"20",x"80",x"00",x"74"),
  1591 => (x"6b",x"63",x"61",x"42"),
  1592 => (x"00",x"12",x"57",x"00"),
  1593 => (x"00",x"2a",x"70",x"00"),
  1594 => (x"00",x"00",x"00",x"00"),
  1595 => (x"00",x"00",x"12",x"57"),
  1596 => (x"00",x"00",x"2a",x"8e"),
  1597 => (x"57",x"00",x"00",x"00"),
  1598 => (x"ac",x"00",x"00",x"12"),
  1599 => (x"00",x"00",x"00",x"2a"),
  1600 => (x"12",x"57",x"00",x"00"),
  1601 => (x"2a",x"ca",x"00",x"00"),
  1602 => (x"00",x"00",x"00",x"00"),
  1603 => (x"00",x"12",x"57",x"00"),
  1604 => (x"00",x"2a",x"e8",x"00"),
  1605 => (x"00",x"00",x"00",x"00"),
  1606 => (x"00",x"00",x"12",x"57"),
  1607 => (x"00",x"00",x"2b",x"06"),
  1608 => (x"57",x"00",x"00",x"00"),
  1609 => (x"24",x"00",x"00",x"12"),
  1610 => (x"00",x"00",x"00",x"2b"),
  1611 => (x"12",x"57",x"00",x"00"),
  1612 => (x"00",x"00",x"00",x"00"),
  1613 => (x"00",x"00",x"00",x"00"),
  1614 => (x"00",x"12",x"ec",x"00"),
  1615 => (x"00",x"00",x"00",x"00"),
  1616 => (x"00",x"00",x"00",x"00"),
  1617 => (x"00",x"00",x"19",x"48"),
  1618 => (x"45",x"53",x"41",x"4c"),
  1619 => (x"30",x"30",x"35",x"52"),
  1620 => (x"00",x"4d",x"4f",x"52"),
  1621 => (x"64",x"61",x"6f",x"4c"),
  1622 => (x"00",x"2e",x"2a",x"20"),
  1623 => (x"48",x"f0",x"fe",x"1e"),
  1624 => (x"09",x"cd",x"78",x"c0"),
  1625 => (x"4f",x"26",x"09",x"79"),
  1626 => (x"f0",x"fe",x"1e",x"1e"),
  1627 => (x"26",x"48",x"7e",x"bf"),
  1628 => (x"fe",x"1e",x"4f",x"26"),
  1629 => (x"78",x"c1",x"48",x"f0"),
  1630 => (x"fe",x"1e",x"4f",x"26"),
  1631 => (x"78",x"c0",x"48",x"f0"),
  1632 => (x"71",x"1e",x"4f",x"26"),
  1633 => (x"52",x"52",x"c0",x"4a"),
  1634 => (x"5e",x"0e",x"4f",x"26"),
  1635 => (x"0e",x"5d",x"5c",x"5b"),
  1636 => (x"4d",x"71",x"86",x"f4"),
  1637 => (x"c1",x"7e",x"6d",x"97"),
  1638 => (x"6c",x"97",x"4c",x"a5"),
  1639 => (x"58",x"a6",x"c8",x"48"),
  1640 => (x"66",x"c4",x"48",x"6e"),
  1641 => (x"87",x"c5",x"05",x"a8"),
  1642 => (x"e6",x"c0",x"48",x"ff"),
  1643 => (x"87",x"ca",x"ff",x"87"),
  1644 => (x"97",x"49",x"a5",x"c2"),
  1645 => (x"a3",x"71",x"4b",x"6c"),
  1646 => (x"4b",x"6b",x"97",x"4b"),
  1647 => (x"6e",x"7e",x"6c",x"97"),
  1648 => (x"c8",x"80",x"c1",x"48"),
  1649 => (x"98",x"c7",x"58",x"a6"),
  1650 => (x"70",x"58",x"a6",x"cc"),
  1651 => (x"e1",x"fe",x"7c",x"97"),
  1652 => (x"f4",x"48",x"73",x"87"),
  1653 => (x"26",x"4d",x"26",x"8e"),
  1654 => (x"26",x"4b",x"26",x"4c"),
  1655 => (x"5b",x"5e",x"0e",x"4f"),
  1656 => (x"86",x"f4",x"0e",x"5c"),
  1657 => (x"66",x"d8",x"4c",x"71"),
  1658 => (x"9a",x"ff",x"c3",x"4a"),
  1659 => (x"97",x"4b",x"a4",x"c2"),
  1660 => (x"a1",x"73",x"49",x"6c"),
  1661 => (x"97",x"51",x"72",x"49"),
  1662 => (x"48",x"6e",x"7e",x"6c"),
  1663 => (x"a6",x"c8",x"80",x"c1"),
  1664 => (x"cc",x"98",x"c7",x"58"),
  1665 => (x"54",x"70",x"58",x"a6"),
  1666 => (x"ca",x"ff",x"8e",x"f4"),
  1667 => (x"fd",x"1e",x"1e",x"87"),
  1668 => (x"bf",x"e0",x"87",x"e8"),
  1669 => (x"e0",x"c0",x"49",x"4a"),
  1670 => (x"cb",x"02",x"99",x"c0"),
  1671 => (x"c2",x"1e",x"72",x"87"),
  1672 => (x"fe",x"49",x"c2",x"ed"),
  1673 => (x"86",x"c4",x"87",x"f7"),
  1674 => (x"70",x"87",x"fd",x"fc"),
  1675 => (x"87",x"c2",x"fd",x"7e"),
  1676 => (x"1e",x"4f",x"26",x"26"),
  1677 => (x"49",x"c2",x"ed",x"c2"),
  1678 => (x"c1",x"87",x"c7",x"fd"),
  1679 => (x"fc",x"49",x"cd",x"e8"),
  1680 => (x"c8",x"c4",x"87",x"da"),
  1681 => (x"1e",x"4f",x"26",x"87"),
  1682 => (x"c8",x"48",x"d0",x"ff"),
  1683 => (x"d4",x"ff",x"78",x"e1"),
  1684 => (x"c4",x"78",x"c5",x"48"),
  1685 => (x"87",x"c3",x"02",x"66"),
  1686 => (x"c8",x"78",x"e0",x"c3"),
  1687 => (x"87",x"c6",x"02",x"66"),
  1688 => (x"c3",x"48",x"d4",x"ff"),
  1689 => (x"d4",x"ff",x"78",x"f0"),
  1690 => (x"ff",x"78",x"71",x"48"),
  1691 => (x"e1",x"c8",x"48",x"d0"),
  1692 => (x"78",x"e0",x"c0",x"78"),
  1693 => (x"5e",x"0e",x"4f",x"26"),
  1694 => (x"71",x"0e",x"5c",x"5b"),
  1695 => (x"c2",x"ed",x"c2",x"4c"),
  1696 => (x"87",x"c6",x"fc",x"49"),
  1697 => (x"b7",x"c0",x"4a",x"70"),
  1698 => (x"e3",x"c2",x"04",x"aa"),
  1699 => (x"aa",x"e0",x"c3",x"87"),
  1700 => (x"c1",x"87",x"c9",x"05"),
  1701 => (x"c1",x"48",x"c0",x"ed"),
  1702 => (x"87",x"d4",x"c2",x"78"),
  1703 => (x"05",x"aa",x"f0",x"c3"),
  1704 => (x"ec",x"c1",x"87",x"c9"),
  1705 => (x"78",x"c1",x"48",x"fc"),
  1706 => (x"c1",x"87",x"f5",x"c1"),
  1707 => (x"02",x"bf",x"c0",x"ed"),
  1708 => (x"4b",x"72",x"87",x"c7"),
  1709 => (x"c2",x"b3",x"c0",x"c2"),
  1710 => (x"74",x"4b",x"72",x"87"),
  1711 => (x"87",x"d1",x"05",x"9c"),
  1712 => (x"bf",x"fc",x"ec",x"c1"),
  1713 => (x"c0",x"ed",x"c1",x"1e"),
  1714 => (x"49",x"72",x"1e",x"bf"),
  1715 => (x"c8",x"87",x"f8",x"fd"),
  1716 => (x"fc",x"ec",x"c1",x"86"),
  1717 => (x"e0",x"c0",x"02",x"bf"),
  1718 => (x"c4",x"49",x"73",x"87"),
  1719 => (x"c1",x"91",x"29",x"b7"),
  1720 => (x"73",x"81",x"dc",x"ee"),
  1721 => (x"c2",x"9a",x"cf",x"4a"),
  1722 => (x"72",x"48",x"c1",x"92"),
  1723 => (x"ff",x"4a",x"70",x"30"),
  1724 => (x"69",x"48",x"72",x"ba"),
  1725 => (x"db",x"79",x"70",x"98"),
  1726 => (x"c4",x"49",x"73",x"87"),
  1727 => (x"c1",x"91",x"29",x"b7"),
  1728 => (x"73",x"81",x"dc",x"ee"),
  1729 => (x"c2",x"9a",x"cf",x"4a"),
  1730 => (x"72",x"48",x"c3",x"92"),
  1731 => (x"48",x"4a",x"70",x"30"),
  1732 => (x"79",x"70",x"b0",x"69"),
  1733 => (x"48",x"c0",x"ed",x"c1"),
  1734 => (x"ec",x"c1",x"78",x"c0"),
  1735 => (x"78",x"c0",x"48",x"fc"),
  1736 => (x"49",x"c2",x"ed",x"c2"),
  1737 => (x"70",x"87",x"e3",x"f9"),
  1738 => (x"aa",x"b7",x"c0",x"4a"),
  1739 => (x"87",x"dd",x"fd",x"03"),
  1740 => (x"87",x"c2",x"48",x"c0"),
  1741 => (x"4c",x"26",x"4d",x"26"),
  1742 => (x"4f",x"26",x"4b",x"26"),
  1743 => (x"00",x"00",x"00",x"00"),
  1744 => (x"00",x"00",x"00",x"00"),
  1745 => (x"49",x"4a",x"71",x"1e"),
  1746 => (x"26",x"87",x"eb",x"fc"),
  1747 => (x"4a",x"c0",x"1e",x"4f"),
  1748 => (x"91",x"c4",x"49",x"72"),
  1749 => (x"81",x"dc",x"ee",x"c1"),
  1750 => (x"82",x"c1",x"79",x"c0"),
  1751 => (x"04",x"aa",x"b7",x"d0"),
  1752 => (x"4f",x"26",x"87",x"ee"),
  1753 => (x"5c",x"5b",x"5e",x"0e"),
  1754 => (x"4d",x"71",x"0e",x"5d"),
  1755 => (x"75",x"87",x"cb",x"f8"),
  1756 => (x"2a",x"b7",x"c4",x"4a"),
  1757 => (x"dc",x"ee",x"c1",x"92"),
  1758 => (x"cf",x"4c",x"75",x"82"),
  1759 => (x"6a",x"94",x"c2",x"9c"),
  1760 => (x"2b",x"74",x"4b",x"49"),
  1761 => (x"48",x"c2",x"9b",x"c3"),
  1762 => (x"4c",x"70",x"30",x"74"),
  1763 => (x"48",x"74",x"bc",x"ff"),
  1764 => (x"7a",x"70",x"98",x"71"),
  1765 => (x"73",x"87",x"db",x"f7"),
  1766 => (x"87",x"d8",x"fe",x"48"),
  1767 => (x"00",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"00",x"00"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"00",x"00",x"00",x"00"),
  1776 => (x"00",x"00",x"00",x"00"),
  1777 => (x"00",x"00",x"00",x"00"),
  1778 => (x"00",x"00",x"00",x"00"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"48",x"d0",x"ff",x"1e"),
  1784 => (x"71",x"78",x"e1",x"c8"),
  1785 => (x"08",x"d4",x"ff",x"48"),
  1786 => (x"1e",x"4f",x"26",x"78"),
  1787 => (x"c8",x"48",x"d0",x"ff"),
  1788 => (x"48",x"71",x"78",x"e1"),
  1789 => (x"78",x"08",x"d4",x"ff"),
  1790 => (x"ff",x"48",x"66",x"c4"),
  1791 => (x"26",x"78",x"08",x"d4"),
  1792 => (x"4a",x"71",x"1e",x"4f"),
  1793 => (x"1e",x"49",x"66",x"c4"),
  1794 => (x"de",x"ff",x"49",x"72"),
  1795 => (x"48",x"d0",x"ff",x"87"),
  1796 => (x"26",x"78",x"e0",x"c0"),
  1797 => (x"73",x"1e",x"4f",x"26"),
  1798 => (x"c8",x"4b",x"71",x"1e"),
  1799 => (x"73",x"1e",x"49",x"66"),
  1800 => (x"a2",x"e0",x"c1",x"4a"),
  1801 => (x"87",x"d9",x"ff",x"49"),
  1802 => (x"26",x"87",x"c4",x"26"),
  1803 => (x"26",x"4c",x"26",x"4d"),
  1804 => (x"1e",x"4f",x"26",x"4b"),
  1805 => (x"c3",x"4a",x"d4",x"ff"),
  1806 => (x"d0",x"ff",x"7a",x"ff"),
  1807 => (x"78",x"e1",x"c8",x"48"),
  1808 => (x"ed",x"c2",x"7a",x"de"),
  1809 => (x"49",x"7a",x"bf",x"cc"),
  1810 => (x"70",x"28",x"c8",x"48"),
  1811 => (x"d0",x"48",x"71",x"7a"),
  1812 => (x"71",x"7a",x"70",x"28"),
  1813 => (x"70",x"28",x"d8",x"48"),
  1814 => (x"48",x"d0",x"ff",x"7a"),
  1815 => (x"26",x"78",x"e0",x"c0"),
  1816 => (x"5b",x"5e",x"0e",x"4f"),
  1817 => (x"71",x"0e",x"5d",x"5c"),
  1818 => (x"cc",x"ed",x"c2",x"4c"),
  1819 => (x"74",x"4b",x"4d",x"bf"),
  1820 => (x"9b",x"66",x"d0",x"2b"),
  1821 => (x"66",x"d4",x"83",x"c1"),
  1822 => (x"87",x"c2",x"04",x"ab"),
  1823 => (x"4a",x"74",x"4b",x"c0"),
  1824 => (x"72",x"49",x"66",x"d0"),
  1825 => (x"75",x"b9",x"ff",x"31"),
  1826 => (x"72",x"48",x"73",x"99"),
  1827 => (x"48",x"4a",x"70",x"30"),
  1828 => (x"ed",x"c2",x"b0",x"71"),
  1829 => (x"da",x"fe",x"58",x"d0"),
  1830 => (x"26",x"4d",x"26",x"87"),
  1831 => (x"26",x"4b",x"26",x"4c"),
  1832 => (x"d0",x"ff",x"1e",x"4f"),
  1833 => (x"78",x"c9",x"c8",x"48"),
  1834 => (x"d4",x"ff",x"48",x"71"),
  1835 => (x"4f",x"26",x"78",x"08"),
  1836 => (x"49",x"4a",x"71",x"1e"),
  1837 => (x"d0",x"ff",x"87",x"eb"),
  1838 => (x"26",x"78",x"c8",x"48"),
  1839 => (x"1e",x"73",x"1e",x"4f"),
  1840 => (x"ed",x"c2",x"4b",x"71"),
  1841 => (x"c3",x"02",x"bf",x"dc"),
  1842 => (x"87",x"eb",x"c2",x"87"),
  1843 => (x"c8",x"48",x"d0",x"ff"),
  1844 => (x"49",x"73",x"78",x"c9"),
  1845 => (x"ff",x"b1",x"e0",x"c0"),
  1846 => (x"78",x"71",x"48",x"d4"),
  1847 => (x"48",x"d0",x"ed",x"c2"),
  1848 => (x"66",x"c8",x"78",x"c0"),
  1849 => (x"c3",x"87",x"c5",x"02"),
  1850 => (x"87",x"c2",x"49",x"ff"),
  1851 => (x"ed",x"c2",x"49",x"c0"),
  1852 => (x"66",x"cc",x"59",x"d8"),
  1853 => (x"c5",x"87",x"c6",x"02"),
  1854 => (x"c4",x"4a",x"d5",x"d5"),
  1855 => (x"ff",x"ff",x"cf",x"87"),
  1856 => (x"dc",x"ed",x"c2",x"4a"),
  1857 => (x"dc",x"ed",x"c2",x"5a"),
  1858 => (x"c4",x"78",x"c1",x"48"),
  1859 => (x"26",x"4d",x"26",x"87"),
  1860 => (x"26",x"4b",x"26",x"4c"),
  1861 => (x"5b",x"5e",x"0e",x"4f"),
  1862 => (x"71",x"0e",x"5d",x"5c"),
  1863 => (x"d8",x"ed",x"c2",x"4a"),
  1864 => (x"9a",x"72",x"4c",x"bf"),
  1865 => (x"49",x"87",x"cb",x"02"),
  1866 => (x"f2",x"c1",x"91",x"c8"),
  1867 => (x"83",x"71",x"4b",x"f3"),
  1868 => (x"f6",x"c1",x"87",x"c4"),
  1869 => (x"4d",x"c0",x"4b",x"f3"),
  1870 => (x"99",x"74",x"49",x"13"),
  1871 => (x"bf",x"d4",x"ed",x"c2"),
  1872 => (x"48",x"d4",x"ff",x"b9"),
  1873 => (x"b7",x"c1",x"78",x"71"),
  1874 => (x"b7",x"c8",x"85",x"2c"),
  1875 => (x"87",x"e8",x"04",x"ad"),
  1876 => (x"bf",x"d0",x"ed",x"c2"),
  1877 => (x"c2",x"80",x"c8",x"48"),
  1878 => (x"fe",x"58",x"d4",x"ed"),
  1879 => (x"73",x"1e",x"87",x"ef"),
  1880 => (x"13",x"4b",x"71",x"1e"),
  1881 => (x"cb",x"02",x"9a",x"4a"),
  1882 => (x"fe",x"49",x"72",x"87"),
  1883 => (x"4a",x"13",x"87",x"e7"),
  1884 => (x"87",x"f5",x"05",x"9a"),
  1885 => (x"1e",x"87",x"da",x"fe"),
  1886 => (x"bf",x"d0",x"ed",x"c2"),
  1887 => (x"d0",x"ed",x"c2",x"49"),
  1888 => (x"78",x"a1",x"c1",x"48"),
  1889 => (x"a9",x"b7",x"c0",x"c4"),
  1890 => (x"ff",x"87",x"db",x"03"),
  1891 => (x"ed",x"c2",x"48",x"d4"),
  1892 => (x"c2",x"78",x"bf",x"d4"),
  1893 => (x"49",x"bf",x"d0",x"ed"),
  1894 => (x"48",x"d0",x"ed",x"c2"),
  1895 => (x"c4",x"78",x"a1",x"c1"),
  1896 => (x"04",x"a9",x"b7",x"c0"),
  1897 => (x"d0",x"ff",x"87",x"e5"),
  1898 => (x"c2",x"78",x"c8",x"48"),
  1899 => (x"c0",x"48",x"dc",x"ed"),
  1900 => (x"00",x"4f",x"26",x"78"),
  1901 => (x"00",x"00",x"00",x"00"),
  1902 => (x"00",x"00",x"00",x"00"),
  1903 => (x"5f",x"5f",x"00",x"00"),
  1904 => (x"00",x"00",x"00",x"00"),
  1905 => (x"03",x"00",x"03",x"03"),
  1906 => (x"14",x"00",x"00",x"03"),
  1907 => (x"7f",x"14",x"7f",x"7f"),
  1908 => (x"00",x"00",x"14",x"7f"),
  1909 => (x"6b",x"6b",x"2e",x"24"),
  1910 => (x"4c",x"00",x"12",x"3a"),
  1911 => (x"6c",x"18",x"36",x"6a"),
  1912 => (x"30",x"00",x"32",x"56"),
  1913 => (x"77",x"59",x"4f",x"7e"),
  1914 => (x"00",x"40",x"68",x"3a"),
  1915 => (x"03",x"07",x"04",x"00"),
  1916 => (x"00",x"00",x"00",x"00"),
  1917 => (x"63",x"3e",x"1c",x"00"),
  1918 => (x"00",x"00",x"00",x"41"),
  1919 => (x"3e",x"63",x"41",x"00"),
  1920 => (x"08",x"00",x"00",x"1c"),
  1921 => (x"1c",x"1c",x"3e",x"2a"),
  1922 => (x"00",x"08",x"2a",x"3e"),
  1923 => (x"3e",x"3e",x"08",x"08"),
  1924 => (x"00",x"00",x"08",x"08"),
  1925 => (x"60",x"e0",x"80",x"00"),
  1926 => (x"00",x"00",x"00",x"00"),
  1927 => (x"08",x"08",x"08",x"08"),
  1928 => (x"00",x"00",x"08",x"08"),
  1929 => (x"60",x"60",x"00",x"00"),
  1930 => (x"40",x"00",x"00",x"00"),
  1931 => (x"0c",x"18",x"30",x"60"),
  1932 => (x"00",x"01",x"03",x"06"),
  1933 => (x"4d",x"59",x"7f",x"3e"),
  1934 => (x"00",x"00",x"3e",x"7f"),
  1935 => (x"7f",x"7f",x"06",x"04"),
  1936 => (x"00",x"00",x"00",x"00"),
  1937 => (x"59",x"71",x"63",x"42"),
  1938 => (x"00",x"00",x"46",x"4f"),
  1939 => (x"49",x"49",x"63",x"22"),
  1940 => (x"18",x"00",x"36",x"7f"),
  1941 => (x"7f",x"13",x"16",x"1c"),
  1942 => (x"00",x"00",x"10",x"7f"),
  1943 => (x"45",x"45",x"67",x"27"),
  1944 => (x"00",x"00",x"39",x"7d"),
  1945 => (x"49",x"4b",x"7e",x"3c"),
  1946 => (x"00",x"00",x"30",x"79"),
  1947 => (x"79",x"71",x"01",x"01"),
  1948 => (x"00",x"00",x"07",x"0f"),
  1949 => (x"49",x"49",x"7f",x"36"),
  1950 => (x"00",x"00",x"36",x"7f"),
  1951 => (x"69",x"49",x"4f",x"06"),
  1952 => (x"00",x"00",x"1e",x"3f"),
  1953 => (x"66",x"66",x"00",x"00"),
  1954 => (x"00",x"00",x"00",x"00"),
  1955 => (x"66",x"e6",x"80",x"00"),
  1956 => (x"00",x"00",x"00",x"00"),
  1957 => (x"14",x"14",x"08",x"08"),
  1958 => (x"00",x"00",x"22",x"22"),
  1959 => (x"14",x"14",x"14",x"14"),
  1960 => (x"00",x"00",x"14",x"14"),
  1961 => (x"14",x"14",x"22",x"22"),
  1962 => (x"00",x"00",x"08",x"08"),
  1963 => (x"59",x"51",x"03",x"02"),
  1964 => (x"3e",x"00",x"06",x"0f"),
  1965 => (x"55",x"5d",x"41",x"7f"),
  1966 => (x"00",x"00",x"1e",x"1f"),
  1967 => (x"09",x"09",x"7f",x"7e"),
  1968 => (x"00",x"00",x"7e",x"7f"),
  1969 => (x"49",x"49",x"7f",x"7f"),
  1970 => (x"00",x"00",x"36",x"7f"),
  1971 => (x"41",x"63",x"3e",x"1c"),
  1972 => (x"00",x"00",x"41",x"41"),
  1973 => (x"63",x"41",x"7f",x"7f"),
  1974 => (x"00",x"00",x"1c",x"3e"),
  1975 => (x"49",x"49",x"7f",x"7f"),
  1976 => (x"00",x"00",x"41",x"41"),
  1977 => (x"09",x"09",x"7f",x"7f"),
  1978 => (x"00",x"00",x"01",x"01"),
  1979 => (x"49",x"41",x"7f",x"3e"),
  1980 => (x"00",x"00",x"7a",x"7b"),
  1981 => (x"08",x"08",x"7f",x"7f"),
  1982 => (x"00",x"00",x"7f",x"7f"),
  1983 => (x"7f",x"7f",x"41",x"00"),
  1984 => (x"00",x"00",x"00",x"41"),
  1985 => (x"40",x"40",x"60",x"20"),
  1986 => (x"7f",x"00",x"3f",x"7f"),
  1987 => (x"36",x"1c",x"08",x"7f"),
  1988 => (x"00",x"00",x"41",x"63"),
  1989 => (x"40",x"40",x"7f",x"7f"),
  1990 => (x"7f",x"00",x"40",x"40"),
  1991 => (x"06",x"0c",x"06",x"7f"),
  1992 => (x"7f",x"00",x"7f",x"7f"),
  1993 => (x"18",x"0c",x"06",x"7f"),
  1994 => (x"00",x"00",x"7f",x"7f"),
  1995 => (x"41",x"41",x"7f",x"3e"),
  1996 => (x"00",x"00",x"3e",x"7f"),
  1997 => (x"09",x"09",x"7f",x"7f"),
  1998 => (x"3e",x"00",x"06",x"0f"),
  1999 => (x"7f",x"61",x"41",x"7f"),
  2000 => (x"00",x"00",x"40",x"7e"),
  2001 => (x"19",x"09",x"7f",x"7f"),
  2002 => (x"00",x"00",x"66",x"7f"),
  2003 => (x"59",x"4d",x"6f",x"26"),
  2004 => (x"00",x"00",x"32",x"7b"),
  2005 => (x"7f",x"7f",x"01",x"01"),
  2006 => (x"00",x"00",x"01",x"01"),
  2007 => (x"40",x"40",x"7f",x"3f"),
  2008 => (x"00",x"00",x"3f",x"7f"),
  2009 => (x"70",x"70",x"3f",x"0f"),
  2010 => (x"7f",x"00",x"0f",x"3f"),
  2011 => (x"30",x"18",x"30",x"7f"),
  2012 => (x"41",x"00",x"7f",x"7f"),
  2013 => (x"1c",x"1c",x"36",x"63"),
  2014 => (x"01",x"41",x"63",x"36"),
  2015 => (x"7c",x"7c",x"06",x"03"),
  2016 => (x"61",x"01",x"03",x"06"),
  2017 => (x"47",x"4d",x"59",x"71"),
  2018 => (x"00",x"00",x"41",x"43"),
  2019 => (x"41",x"7f",x"7f",x"00"),
  2020 => (x"01",x"00",x"00",x"41"),
  2021 => (x"18",x"0c",x"06",x"03"),
  2022 => (x"00",x"40",x"60",x"30"),
  2023 => (x"7f",x"41",x"41",x"00"),
  2024 => (x"08",x"00",x"00",x"7f"),
  2025 => (x"06",x"03",x"06",x"0c"),
  2026 => (x"80",x"00",x"08",x"0c"),
  2027 => (x"80",x"80",x"80",x"80"),
  2028 => (x"00",x"00",x"80",x"80"),
  2029 => (x"07",x"03",x"00",x"00"),
  2030 => (x"00",x"00",x"00",x"04"),
  2031 => (x"54",x"54",x"74",x"20"),
  2032 => (x"00",x"00",x"78",x"7c"),
  2033 => (x"44",x"44",x"7f",x"7f"),
  2034 => (x"00",x"00",x"38",x"7c"),
  2035 => (x"44",x"44",x"7c",x"38"),
  2036 => (x"00",x"00",x"00",x"44"),
  2037 => (x"44",x"44",x"7c",x"38"),
  2038 => (x"00",x"00",x"7f",x"7f"),
  2039 => (x"54",x"54",x"7c",x"38"),
  2040 => (x"00",x"00",x"18",x"5c"),
  2041 => (x"05",x"7f",x"7e",x"04"),
  2042 => (x"00",x"00",x"00",x"05"),
  2043 => (x"a4",x"a4",x"bc",x"18"),
  2044 => (x"00",x"00",x"7c",x"fc"),
  2045 => (x"04",x"04",x"7f",x"7f"),
  2046 => (x"00",x"00",x"78",x"7c"),
  2047 => (x"7d",x"3d",x"00",x"00"),
  2048 => (x"00",x"00",x"00",x"40"),
  2049 => (x"fd",x"80",x"80",x"80"),
  2050 => (x"00",x"00",x"00",x"7d"),
  2051 => (x"38",x"10",x"7f",x"7f"),
  2052 => (x"00",x"00",x"44",x"6c"),
  2053 => (x"7f",x"3f",x"00",x"00"),
  2054 => (x"7c",x"00",x"00",x"40"),
  2055 => (x"0c",x"18",x"0c",x"7c"),
  2056 => (x"00",x"00",x"78",x"7c"),
  2057 => (x"04",x"04",x"7c",x"7c"),
  2058 => (x"00",x"00",x"78",x"7c"),
  2059 => (x"44",x"44",x"7c",x"38"),
  2060 => (x"00",x"00",x"38",x"7c"),
  2061 => (x"24",x"24",x"fc",x"fc"),
  2062 => (x"00",x"00",x"18",x"3c"),
  2063 => (x"24",x"24",x"3c",x"18"),
  2064 => (x"00",x"00",x"fc",x"fc"),
  2065 => (x"04",x"04",x"7c",x"7c"),
  2066 => (x"00",x"00",x"08",x"0c"),
  2067 => (x"54",x"54",x"5c",x"48"),
  2068 => (x"00",x"00",x"20",x"74"),
  2069 => (x"44",x"7f",x"3f",x"04"),
  2070 => (x"00",x"00",x"00",x"44"),
  2071 => (x"40",x"40",x"7c",x"3c"),
  2072 => (x"00",x"00",x"7c",x"7c"),
  2073 => (x"60",x"60",x"3c",x"1c"),
  2074 => (x"3c",x"00",x"1c",x"3c"),
  2075 => (x"60",x"30",x"60",x"7c"),
  2076 => (x"44",x"00",x"3c",x"7c"),
  2077 => (x"38",x"10",x"38",x"6c"),
  2078 => (x"00",x"00",x"44",x"6c"),
  2079 => (x"60",x"e0",x"bc",x"1c"),
  2080 => (x"00",x"00",x"1c",x"3c"),
  2081 => (x"5c",x"74",x"64",x"44"),
  2082 => (x"00",x"00",x"44",x"4c"),
  2083 => (x"77",x"3e",x"08",x"08"),
  2084 => (x"00",x"00",x"41",x"41"),
  2085 => (x"7f",x"7f",x"00",x"00"),
  2086 => (x"00",x"00",x"00",x"00"),
  2087 => (x"3e",x"77",x"41",x"41"),
  2088 => (x"02",x"00",x"08",x"08"),
  2089 => (x"02",x"03",x"01",x"01"),
  2090 => (x"7f",x"00",x"01",x"02"),
  2091 => (x"7f",x"7f",x"7f",x"7f"),
  2092 => (x"08",x"00",x"7f",x"7f"),
  2093 => (x"3e",x"1c",x"1c",x"08"),
  2094 => (x"7f",x"7f",x"7f",x"3e"),
  2095 => (x"1c",x"3e",x"3e",x"7f"),
  2096 => (x"00",x"08",x"08",x"1c"),
  2097 => (x"7c",x"7c",x"18",x"10"),
  2098 => (x"00",x"00",x"10",x"18"),
  2099 => (x"7c",x"7c",x"30",x"10"),
  2100 => (x"10",x"00",x"10",x"30"),
  2101 => (x"78",x"60",x"60",x"30"),
  2102 => (x"42",x"00",x"06",x"1e"),
  2103 => (x"3c",x"18",x"3c",x"66"),
  2104 => (x"78",x"00",x"42",x"66"),
  2105 => (x"c6",x"c2",x"6a",x"38"),
  2106 => (x"60",x"00",x"38",x"6c"),
  2107 => (x"00",x"60",x"00",x"00"),
  2108 => (x"0e",x"00",x"60",x"00"),
  2109 => (x"5d",x"5c",x"5b",x"5e"),
  2110 => (x"4c",x"71",x"1e",x"0e"),
  2111 => (x"bf",x"ed",x"ed",x"c2"),
  2112 => (x"c0",x"4b",x"c0",x"4d"),
  2113 => (x"02",x"ab",x"74",x"1e"),
  2114 => (x"a6",x"c4",x"87",x"c7"),
  2115 => (x"c5",x"78",x"c0",x"48"),
  2116 => (x"48",x"a6",x"c4",x"87"),
  2117 => (x"66",x"c4",x"78",x"c1"),
  2118 => (x"ee",x"49",x"73",x"1e"),
  2119 => (x"86",x"c8",x"87",x"df"),
  2120 => (x"ef",x"49",x"e0",x"c0"),
  2121 => (x"a5",x"c4",x"87",x"ef"),
  2122 => (x"f0",x"49",x"6a",x"4a"),
  2123 => (x"c6",x"f1",x"87",x"f0"),
  2124 => (x"c1",x"85",x"cb",x"87"),
  2125 => (x"ab",x"b7",x"c8",x"83"),
  2126 => (x"87",x"c7",x"ff",x"04"),
  2127 => (x"26",x"4d",x"26",x"26"),
  2128 => (x"26",x"4b",x"26",x"4c"),
  2129 => (x"4a",x"71",x"1e",x"4f"),
  2130 => (x"5a",x"f1",x"ed",x"c2"),
  2131 => (x"48",x"f1",x"ed",x"c2"),
  2132 => (x"fe",x"49",x"78",x"c7"),
  2133 => (x"4f",x"26",x"87",x"dd"),
  2134 => (x"71",x"1e",x"73",x"1e"),
  2135 => (x"aa",x"b7",x"c0",x"4a"),
  2136 => (x"c2",x"87",x"d3",x"03"),
  2137 => (x"05",x"bf",x"e8",x"d2"),
  2138 => (x"4b",x"c1",x"87",x"c4"),
  2139 => (x"4b",x"c0",x"87",x"c2"),
  2140 => (x"5b",x"ec",x"d2",x"c2"),
  2141 => (x"d2",x"c2",x"87",x"c4"),
  2142 => (x"d2",x"c2",x"5a",x"ec"),
  2143 => (x"c1",x"4a",x"bf",x"e8"),
  2144 => (x"a2",x"c0",x"c1",x"9a"),
  2145 => (x"87",x"e8",x"ec",x"49"),
  2146 => (x"d2",x"c2",x"48",x"fc"),
  2147 => (x"fe",x"78",x"bf",x"e8"),
  2148 => (x"71",x"1e",x"87",x"ef"),
  2149 => (x"1e",x"66",x"c4",x"4a"),
  2150 => (x"f9",x"e9",x"49",x"72"),
  2151 => (x"4f",x"26",x"26",x"87"),
  2152 => (x"e8",x"d2",x"c2",x"1e"),
  2153 => (x"db",x"e6",x"49",x"bf"),
  2154 => (x"e5",x"ed",x"c2",x"87"),
  2155 => (x"78",x"bf",x"e8",x"48"),
  2156 => (x"48",x"e1",x"ed",x"c2"),
  2157 => (x"c2",x"78",x"bf",x"ec"),
  2158 => (x"4a",x"bf",x"e5",x"ed"),
  2159 => (x"99",x"ff",x"c3",x"49"),
  2160 => (x"72",x"2a",x"b7",x"c8"),
  2161 => (x"c2",x"b0",x"71",x"48"),
  2162 => (x"26",x"58",x"ed",x"ed"),
  2163 => (x"5b",x"5e",x"0e",x"4f"),
  2164 => (x"71",x"0e",x"5d",x"5c"),
  2165 => (x"87",x"c8",x"ff",x"4b"),
  2166 => (x"48",x"e0",x"ed",x"c2"),
  2167 => (x"49",x"73",x"50",x"c0"),
  2168 => (x"70",x"87",x"c1",x"e6"),
  2169 => (x"9c",x"c2",x"4c",x"49"),
  2170 => (x"cb",x"49",x"ee",x"cb"),
  2171 => (x"49",x"70",x"87",x"c2"),
  2172 => (x"e0",x"ed",x"c2",x"4d"),
  2173 => (x"c1",x"05",x"bf",x"97"),
  2174 => (x"66",x"d0",x"87",x"e2"),
  2175 => (x"e9",x"ed",x"c2",x"49"),
  2176 => (x"d6",x"05",x"99",x"bf"),
  2177 => (x"49",x"66",x"d4",x"87"),
  2178 => (x"bf",x"e1",x"ed",x"c2"),
  2179 => (x"87",x"cb",x"05",x"99"),
  2180 => (x"cf",x"e5",x"49",x"73"),
  2181 => (x"02",x"98",x"70",x"87"),
  2182 => (x"c1",x"87",x"c1",x"c1"),
  2183 => (x"87",x"c0",x"fe",x"4c"),
  2184 => (x"d7",x"ca",x"49",x"75"),
  2185 => (x"02",x"98",x"70",x"87"),
  2186 => (x"ed",x"c2",x"87",x"c6"),
  2187 => (x"50",x"c1",x"48",x"e0"),
  2188 => (x"97",x"e0",x"ed",x"c2"),
  2189 => (x"e3",x"c0",x"05",x"bf"),
  2190 => (x"e9",x"ed",x"c2",x"87"),
  2191 => (x"66",x"d0",x"49",x"bf"),
  2192 => (x"d6",x"ff",x"05",x"99"),
  2193 => (x"e1",x"ed",x"c2",x"87"),
  2194 => (x"66",x"d4",x"49",x"bf"),
  2195 => (x"ca",x"ff",x"05",x"99"),
  2196 => (x"e4",x"49",x"73",x"87"),
  2197 => (x"98",x"70",x"87",x"ce"),
  2198 => (x"87",x"ff",x"fe",x"05"),
  2199 => (x"dc",x"fb",x"48",x"74"),
  2200 => (x"5b",x"5e",x"0e",x"87"),
  2201 => (x"f4",x"0e",x"5d",x"5c"),
  2202 => (x"4c",x"4d",x"c0",x"86"),
  2203 => (x"c4",x"7e",x"bf",x"ec"),
  2204 => (x"ed",x"c2",x"48",x"a6"),
  2205 => (x"c1",x"78",x"bf",x"ed"),
  2206 => (x"c7",x"1e",x"c0",x"1e"),
  2207 => (x"87",x"cd",x"fd",x"49"),
  2208 => (x"98",x"70",x"86",x"c8"),
  2209 => (x"ff",x"87",x"cd",x"02"),
  2210 => (x"87",x"cc",x"fb",x"49"),
  2211 => (x"e3",x"49",x"da",x"c1"),
  2212 => (x"4d",x"c1",x"87",x"d2"),
  2213 => (x"97",x"e0",x"ed",x"c2"),
  2214 => (x"87",x"c3",x"02",x"bf"),
  2215 => (x"c2",x"87",x"fb",x"cf"),
  2216 => (x"4b",x"bf",x"e5",x"ed"),
  2217 => (x"bf",x"e8",x"d2",x"c2"),
  2218 => (x"87",x"e9",x"c0",x"05"),
  2219 => (x"e2",x"49",x"fd",x"c3"),
  2220 => (x"fa",x"c3",x"87",x"f2"),
  2221 => (x"87",x"ec",x"e2",x"49"),
  2222 => (x"ff",x"c3",x"49",x"73"),
  2223 => (x"c0",x"1e",x"71",x"99"),
  2224 => (x"87",x"ce",x"fb",x"49"),
  2225 => (x"b7",x"c8",x"49",x"73"),
  2226 => (x"c1",x"1e",x"71",x"29"),
  2227 => (x"87",x"c2",x"fb",x"49"),
  2228 => (x"f9",x"c5",x"86",x"c8"),
  2229 => (x"e9",x"ed",x"c2",x"87"),
  2230 => (x"02",x"9b",x"4b",x"bf"),
  2231 => (x"d2",x"c2",x"87",x"dd"),
  2232 => (x"c7",x"49",x"bf",x"e4"),
  2233 => (x"98",x"70",x"87",x"d6"),
  2234 => (x"c0",x"87",x"c4",x"05"),
  2235 => (x"c2",x"87",x"d2",x"4b"),
  2236 => (x"fb",x"c6",x"49",x"e0"),
  2237 => (x"e8",x"d2",x"c2",x"87"),
  2238 => (x"c2",x"87",x"c6",x"58"),
  2239 => (x"c0",x"48",x"e4",x"d2"),
  2240 => (x"c2",x"49",x"73",x"78"),
  2241 => (x"87",x"cd",x"05",x"99"),
  2242 => (x"e1",x"49",x"eb",x"c3"),
  2243 => (x"49",x"70",x"87",x"d6"),
  2244 => (x"c2",x"02",x"99",x"c2"),
  2245 => (x"73",x"4c",x"fb",x"87"),
  2246 => (x"05",x"99",x"c1",x"49"),
  2247 => (x"f4",x"c3",x"87",x"cd"),
  2248 => (x"87",x"c0",x"e1",x"49"),
  2249 => (x"99",x"c2",x"49",x"70"),
  2250 => (x"fa",x"87",x"c2",x"02"),
  2251 => (x"c8",x"49",x"73",x"4c"),
  2252 => (x"87",x"cd",x"05",x"99"),
  2253 => (x"e0",x"49",x"f5",x"c3"),
  2254 => (x"49",x"70",x"87",x"ea"),
  2255 => (x"d4",x"02",x"99",x"c2"),
  2256 => (x"f1",x"ed",x"c2",x"87"),
  2257 => (x"87",x"c9",x"02",x"bf"),
  2258 => (x"c2",x"88",x"c1",x"48"),
  2259 => (x"c2",x"58",x"f5",x"ed"),
  2260 => (x"c1",x"4c",x"ff",x"87"),
  2261 => (x"c4",x"49",x"73",x"4d"),
  2262 => (x"87",x"cd",x"05",x"99"),
  2263 => (x"e0",x"49",x"f2",x"c3"),
  2264 => (x"49",x"70",x"87",x"c2"),
  2265 => (x"db",x"02",x"99",x"c2"),
  2266 => (x"f1",x"ed",x"c2",x"87"),
  2267 => (x"c7",x"48",x"7e",x"bf"),
  2268 => (x"cb",x"03",x"a8",x"b7"),
  2269 => (x"c1",x"48",x"6e",x"87"),
  2270 => (x"f5",x"ed",x"c2",x"80"),
  2271 => (x"87",x"c2",x"c0",x"58"),
  2272 => (x"4d",x"c1",x"4c",x"fe"),
  2273 => (x"ff",x"49",x"fd",x"c3"),
  2274 => (x"70",x"87",x"d9",x"df"),
  2275 => (x"02",x"99",x"c2",x"49"),
  2276 => (x"ed",x"c2",x"87",x"d5"),
  2277 => (x"c0",x"02",x"bf",x"f1"),
  2278 => (x"ed",x"c2",x"87",x"c9"),
  2279 => (x"78",x"c0",x"48",x"f1"),
  2280 => (x"fd",x"87",x"c2",x"c0"),
  2281 => (x"c3",x"4d",x"c1",x"4c"),
  2282 => (x"de",x"ff",x"49",x"fa"),
  2283 => (x"49",x"70",x"87",x"f6"),
  2284 => (x"d9",x"02",x"99",x"c2"),
  2285 => (x"f1",x"ed",x"c2",x"87"),
  2286 => (x"b7",x"c7",x"48",x"bf"),
  2287 => (x"c9",x"c0",x"03",x"a8"),
  2288 => (x"f1",x"ed",x"c2",x"87"),
  2289 => (x"c0",x"78",x"c7",x"48"),
  2290 => (x"4c",x"fc",x"87",x"c2"),
  2291 => (x"b7",x"c0",x"4d",x"c1"),
  2292 => (x"d1",x"c0",x"03",x"ac"),
  2293 => (x"4a",x"66",x"c4",x"87"),
  2294 => (x"6a",x"82",x"d8",x"c1"),
  2295 => (x"87",x"c6",x"c0",x"02"),
  2296 => (x"49",x"74",x"4b",x"6a"),
  2297 => (x"1e",x"c0",x"0f",x"73"),
  2298 => (x"c1",x"1e",x"f0",x"c3"),
  2299 => (x"dc",x"f7",x"49",x"da"),
  2300 => (x"70",x"86",x"c8",x"87"),
  2301 => (x"e2",x"c0",x"02",x"98"),
  2302 => (x"48",x"a6",x"c8",x"87"),
  2303 => (x"bf",x"f1",x"ed",x"c2"),
  2304 => (x"49",x"66",x"c8",x"78"),
  2305 => (x"66",x"c4",x"91",x"cb"),
  2306 => (x"70",x"80",x"71",x"48"),
  2307 => (x"02",x"bf",x"6e",x"7e"),
  2308 => (x"6e",x"87",x"c8",x"c0"),
  2309 => (x"66",x"c8",x"4b",x"bf"),
  2310 => (x"75",x"0f",x"73",x"49"),
  2311 => (x"c8",x"c0",x"02",x"9d"),
  2312 => (x"f1",x"ed",x"c2",x"87"),
  2313 => (x"ca",x"f3",x"49",x"bf"),
  2314 => (x"ec",x"d2",x"c2",x"87"),
  2315 => (x"dd",x"c0",x"02",x"bf"),
  2316 => (x"c7",x"c2",x"49",x"87"),
  2317 => (x"02",x"98",x"70",x"87"),
  2318 => (x"c2",x"87",x"d3",x"c0"),
  2319 => (x"49",x"bf",x"f1",x"ed"),
  2320 => (x"c0",x"87",x"f0",x"f2"),
  2321 => (x"87",x"d0",x"f4",x"49"),
  2322 => (x"48",x"ec",x"d2",x"c2"),
  2323 => (x"8e",x"f4",x"78",x"c0"),
  2324 => (x"0e",x"87",x"ea",x"f3"),
  2325 => (x"5d",x"5c",x"5b",x"5e"),
  2326 => (x"4c",x"71",x"1e",x"0e"),
  2327 => (x"bf",x"ed",x"ed",x"c2"),
  2328 => (x"a1",x"cd",x"c1",x"49"),
  2329 => (x"81",x"d1",x"c1",x"4d"),
  2330 => (x"9c",x"74",x"7e",x"69"),
  2331 => (x"c4",x"87",x"cf",x"02"),
  2332 => (x"7b",x"74",x"4b",x"a5"),
  2333 => (x"bf",x"ed",x"ed",x"c2"),
  2334 => (x"87",x"c9",x"f3",x"49"),
  2335 => (x"9c",x"74",x"7b",x"6e"),
  2336 => (x"c0",x"87",x"c4",x"05"),
  2337 => (x"c1",x"87",x"c2",x"4b"),
  2338 => (x"f3",x"49",x"73",x"4b"),
  2339 => (x"66",x"d4",x"87",x"ca"),
  2340 => (x"49",x"87",x"c7",x"02"),
  2341 => (x"4a",x"70",x"87",x"da"),
  2342 => (x"4a",x"c0",x"87",x"c2"),
  2343 => (x"5a",x"f0",x"d2",x"c2"),
  2344 => (x"87",x"d9",x"f2",x"26"),
  2345 => (x"00",x"00",x"00",x"00"),
  2346 => (x"00",x"00",x"00",x"00"),
  2347 => (x"00",x"00",x"00",x"00"),
  2348 => (x"ff",x"4a",x"71",x"1e"),
  2349 => (x"72",x"49",x"bf",x"c8"),
  2350 => (x"4f",x"26",x"48",x"a1"),
  2351 => (x"bf",x"c8",x"ff",x"1e"),
  2352 => (x"c0",x"c0",x"fe",x"89"),
  2353 => (x"a9",x"c0",x"c0",x"c0"),
  2354 => (x"c0",x"87",x"c4",x"01"),
  2355 => (x"c1",x"87",x"c2",x"4a"),
  2356 => (x"26",x"48",x"72",x"4a"),
  2357 => (x"5b",x"5e",x"0e",x"4f"),
  2358 => (x"71",x"0e",x"5d",x"5c"),
  2359 => (x"4c",x"d4",x"ff",x"4b"),
  2360 => (x"c0",x"48",x"66",x"d0"),
  2361 => (x"ff",x"49",x"d6",x"78"),
  2362 => (x"c3",x"87",x"f1",x"db"),
  2363 => (x"49",x"6c",x"7c",x"ff"),
  2364 => (x"71",x"99",x"ff",x"c3"),
  2365 => (x"f0",x"c3",x"49",x"4d"),
  2366 => (x"a9",x"e0",x"c1",x"99"),
  2367 => (x"c3",x"87",x"cb",x"05"),
  2368 => (x"48",x"6c",x"7c",x"ff"),
  2369 => (x"66",x"d0",x"98",x"c3"),
  2370 => (x"ff",x"c3",x"78",x"08"),
  2371 => (x"49",x"4a",x"6c",x"7c"),
  2372 => (x"ff",x"c3",x"31",x"c8"),
  2373 => (x"71",x"4a",x"6c",x"7c"),
  2374 => (x"c8",x"49",x"72",x"b2"),
  2375 => (x"7c",x"ff",x"c3",x"31"),
  2376 => (x"b2",x"71",x"4a",x"6c"),
  2377 => (x"31",x"c8",x"49",x"72"),
  2378 => (x"6c",x"7c",x"ff",x"c3"),
  2379 => (x"ff",x"b2",x"71",x"4a"),
  2380 => (x"e0",x"c0",x"48",x"d0"),
  2381 => (x"02",x"9b",x"73",x"78"),
  2382 => (x"7b",x"72",x"87",x"c2"),
  2383 => (x"4d",x"26",x"48",x"75"),
  2384 => (x"4b",x"26",x"4c",x"26"),
  2385 => (x"26",x"1e",x"4f",x"26"),
  2386 => (x"5b",x"5e",x"0e",x"4f"),
  2387 => (x"86",x"f8",x"0e",x"5c"),
  2388 => (x"a6",x"c8",x"1e",x"76"),
  2389 => (x"87",x"fd",x"fd",x"49"),
  2390 => (x"4b",x"70",x"86",x"c4"),
  2391 => (x"a8",x"c2",x"48",x"6e"),
  2392 => (x"87",x"f0",x"c2",x"03"),
  2393 => (x"f0",x"c3",x"4a",x"73"),
  2394 => (x"aa",x"d0",x"c1",x"9a"),
  2395 => (x"c1",x"87",x"c7",x"02"),
  2396 => (x"c2",x"05",x"aa",x"e0"),
  2397 => (x"49",x"73",x"87",x"de"),
  2398 => (x"c3",x"02",x"99",x"c8"),
  2399 => (x"87",x"c6",x"ff",x"87"),
  2400 => (x"9c",x"c3",x"4c",x"73"),
  2401 => (x"c1",x"05",x"ac",x"c2"),
  2402 => (x"66",x"c4",x"87",x"c2"),
  2403 => (x"71",x"31",x"c9",x"49"),
  2404 => (x"4a",x"66",x"c4",x"1e"),
  2405 => (x"ed",x"c2",x"92",x"d4"),
  2406 => (x"81",x"72",x"49",x"f5"),
  2407 => (x"87",x"c0",x"d1",x"fe"),
  2408 => (x"d8",x"ff",x"49",x"d8"),
  2409 => (x"c0",x"c8",x"87",x"f6"),
  2410 => (x"d2",x"dc",x"c2",x"1e"),
  2411 => (x"fb",x"ec",x"fd",x"49"),
  2412 => (x"48",x"d0",x"ff",x"87"),
  2413 => (x"c2",x"78",x"e0",x"c0"),
  2414 => (x"cc",x"1e",x"d2",x"dc"),
  2415 => (x"92",x"d4",x"4a",x"66"),
  2416 => (x"49",x"f5",x"ed",x"c2"),
  2417 => (x"cf",x"fe",x"81",x"72"),
  2418 => (x"86",x"cc",x"87",x"c7"),
  2419 => (x"c1",x"05",x"ac",x"c1"),
  2420 => (x"66",x"c4",x"87",x"c2"),
  2421 => (x"71",x"31",x"c9",x"49"),
  2422 => (x"4a",x"66",x"c4",x"1e"),
  2423 => (x"ed",x"c2",x"92",x"d4"),
  2424 => (x"81",x"72",x"49",x"f5"),
  2425 => (x"87",x"f8",x"cf",x"fe"),
  2426 => (x"1e",x"d2",x"dc",x"c2"),
  2427 => (x"d4",x"4a",x"66",x"c8"),
  2428 => (x"f5",x"ed",x"c2",x"92"),
  2429 => (x"fe",x"81",x"72",x"49"),
  2430 => (x"d7",x"87",x"c7",x"cd"),
  2431 => (x"db",x"d7",x"ff",x"49"),
  2432 => (x"1e",x"c0",x"c8",x"87"),
  2433 => (x"49",x"d2",x"dc",x"c2"),
  2434 => (x"87",x"f9",x"ea",x"fd"),
  2435 => (x"d0",x"ff",x"86",x"cc"),
  2436 => (x"78",x"e0",x"c0",x"48"),
  2437 => (x"e7",x"fc",x"8e",x"f8"),
  2438 => (x"5b",x"5e",x"0e",x"87"),
  2439 => (x"1e",x"0e",x"5d",x"5c"),
  2440 => (x"d4",x"ff",x"4d",x"71"),
  2441 => (x"7e",x"66",x"d4",x"4c"),
  2442 => (x"a8",x"b7",x"c3",x"48"),
  2443 => (x"c0",x"87",x"c5",x"06"),
  2444 => (x"87",x"e2",x"c1",x"48"),
  2445 => (x"dd",x"fe",x"49",x"75"),
  2446 => (x"1e",x"75",x"87",x"fb"),
  2447 => (x"d4",x"4b",x"66",x"c4"),
  2448 => (x"f5",x"ed",x"c2",x"93"),
  2449 => (x"fe",x"49",x"73",x"83"),
  2450 => (x"c8",x"87",x"e2",x"c8"),
  2451 => (x"ff",x"4b",x"6b",x"83"),
  2452 => (x"e1",x"c8",x"48",x"d0"),
  2453 => (x"73",x"7c",x"dd",x"78"),
  2454 => (x"99",x"ff",x"c3",x"49"),
  2455 => (x"49",x"73",x"7c",x"71"),
  2456 => (x"c3",x"29",x"b7",x"c8"),
  2457 => (x"7c",x"71",x"99",x"ff"),
  2458 => (x"b7",x"d0",x"49",x"73"),
  2459 => (x"99",x"ff",x"c3",x"29"),
  2460 => (x"49",x"73",x"7c",x"71"),
  2461 => (x"71",x"29",x"b7",x"d8"),
  2462 => (x"7c",x"7c",x"c0",x"7c"),
  2463 => (x"7c",x"7c",x"7c",x"7c"),
  2464 => (x"7c",x"7c",x"7c",x"7c"),
  2465 => (x"e0",x"c0",x"7c",x"7c"),
  2466 => (x"1e",x"66",x"c4",x"78"),
  2467 => (x"d5",x"ff",x"49",x"dc"),
  2468 => (x"86",x"c8",x"87",x"ef"),
  2469 => (x"fa",x"26",x"48",x"73"),
  2470 => (x"c2",x"1e",x"87",x"e4"),
  2471 => (x"49",x"bf",x"e8",x"db"),
  2472 => (x"db",x"c2",x"b9",x"c1"),
  2473 => (x"d4",x"ff",x"59",x"ec"),
  2474 => (x"78",x"ff",x"c3",x"48"),
  2475 => (x"c8",x"48",x"d0",x"ff"),
  2476 => (x"d4",x"ff",x"78",x"e1"),
  2477 => (x"c4",x"78",x"c1",x"48"),
  2478 => (x"ff",x"78",x"71",x"31"),
  2479 => (x"e0",x"c0",x"48",x"d0"),
  2480 => (x"1e",x"4f",x"26",x"78"),
  2481 => (x"1e",x"dc",x"db",x"c2"),
  2482 => (x"49",x"c8",x"e9",x"c2"),
  2483 => (x"87",x"dd",x"c6",x"fe"),
  2484 => (x"98",x"70",x"86",x"c4"),
  2485 => (x"ff",x"87",x"c3",x"02"),
  2486 => (x"4f",x"26",x"87",x"c0"),
  2487 => (x"48",x"4b",x"35",x"31"),
  2488 => (x"20",x"20",x"20",x"5a"),
  2489 => (x"00",x"47",x"46",x"43"),
  2490 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

